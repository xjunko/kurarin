module dummy

// Dummy audio backend - might no need this.
fn init() {}
