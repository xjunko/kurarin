module beatmap

import framework.math.time

import object
import timing

// god i fucking hate typescript/javascript
// source: https://github.com/NonSpicyBurrito/sonolus-pjsekai-engine/blob/d2a3c6bda1ef43502e77dcc39cb6e965f86cec7e/src/lib/sus/analyze.ts#L3

pub const (
		ticks_per_beat = 480.0
		ticks_per_hidden = ticks_per_beat / 2.0
)

// Structs
pub struct Line {
	pub mut:
		header string
		data string
}

pub struct MeasureChange {
	pub mut:
		a f64
		b f64
}

pub struct BarLength {
	pub mut:
		measure f64
		length f64
}

pub struct Bar {
	pub mut:
		measure f64
		ticks_per_measure f64
		ticks f64
}

pub struct RawObject {
	pub mut:
		tick f64
		value string
}
//

pub struct Beatmap {
	pub mut:
		lines   []Line
		measure []MeasureChange
		bars []Bar
		barlengths []BarLength
		meta    map[string]string
		
		bpms map[string]f64
		bpm_changes []RawObject
		tap_notes []object.NoteObject
		directional_notes []object.NoteObject
		stream map[string]object.NoteObject

		timings timing.Timing
}

// Resolver
pub fn (mut beatmap Beatmap) resolve_object_time() {
	for mut note in beatmap.tap_notes {
		time := beatmap.to_time(note.tick)
		note.time.start = time
		note.time.end = time
	}
}

pub fn (mut beatmap Beatmap) resolve_note_sprite() {

}

// Time converters
pub fn (mut beatmap Beatmap) to_tick(measure f64, p f64, q f64) f64 {
	mut bar := Bar{ticks: 0xDEAD}

	for bar_to_find in beatmap.bars {
		if measure >= bar_to_find.measure {
			bar = bar_to_find
			break
		}
	}

	if bar.ticks == 0xDEAD { panic("Invalid bar") }

	return bar.ticks + 
		(measure - bar.measure) * bar.ticks_per_measure +
		(p * bar.ticks_per_measure) / q
}

pub fn (mut beatmap Beatmap) to_time(tick f64) f64 {
	return beatmap.timings.to_time(tick)
}