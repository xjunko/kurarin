module object
