module constants

pub const game_name = 'Kurarin'
pub const game_version = 'rewrite-0.0.6.5 [osu!]'
