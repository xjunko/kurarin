module ruleset

pub enum HitResult {
	ignore
	slider_miss
	miss
	hit50
	hit100
	hit300
}