module elzma

pub fn decode_lzma(data []u8) !string {
	return ''
}
