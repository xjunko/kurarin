module object

import framework.math.time

pub struct BaseNoteObject {
	pub mut:
		time time.Time
}