module sekai

import core.sekai.beatmap

import framework.logging

pub fn main() {
	logging.error("${@MOD}: game loop not done yet.")
}