module constants

pub const (
	game_name = "Kurarin"
	game_version = "rewrite-0.0.2b-preview-gui1"
)