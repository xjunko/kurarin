module context

pub fn vsync(enable bool) {
}
