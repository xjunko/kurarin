module sprite

/*
import gx

import framework.math.vector

// will not be used until v support embedded struct on interface
pub struct TextSprite {
	Sprite

	pub mut:
		text string
}

pub fn (s TextSprite) add_transform(arg AddTransformArgument) {

}

pub fn (s TextSprite) after_add_transform_reset() {

}

pub fn (s TextSprite) change_size(t vector.Vector2) {

}


pub fn (s TextSprite) draw(cfg DrawConfig) {
	/*
	if !s.check_if_drawable(cfg.time) && !s.always_visible { return }

	mut img := s.image()

	x := int((s.position.x * cfg.scale - (s.size.x * cfg.scale) / 2) + cfg.offset.x * cfg.scale)
	y := int((s.position.y * cfg.scale - (s.size.x * cfg.scale) / 2) + cfg.offset.y * cfg.scale)
	width := int(s.size.x * cfg.scale)

	cfg.ctx.draw_text(x, y, s.text, gx.TextCfg{
		color: s.color,
		size: width,
		align: .center
	})
	*/
}	

pub fn (s TextSprite) draw_and_update(cfg DrawConfig) {
	/*
	if !s.check_if_drawable(cfg.time) && !s.always_visible { return }

	mut img := s.image()

	x := int((s.position.x * cfg.scale - (s.size.x * cfg.scale) / 2) + cfg.offset.x * cfg.scale)
	y := int((s.position.y * cfg.scale - (s.size.x * cfg.scale) / 2) + cfg.offset.y * cfg.scale)
	width := int(s.size.x * cfg.scale)

	cfg.ctx.draw_text(x, y, s.text, gx.TextCfg{
		color: s.color,
		size: width,
		align: .center
	})
	*/
}	

*/