module cursor

import math

import game.beatmap
import game.beatmap.object as gameobject
import game.movers

import framework.math.time
import framework.math.vector
import framework.math.easing

import game.settings

const (
	offset = settings.gameplay.auto_update_rate
)

[deprecated: "TODO: remove this after we got realtime auto."]
pub fn make_replay(mut beatmap &beatmap.Beatmap, mut cursor &Cursor) {
	mut last_object := unsafe { &beatmap.objects[0] }
	mut last_position := beatmap.objects[0].get_start_position()
	mut direction := 1

	for mut object in beatmap.objects {
		if mut object is gameobject.Circle || mut object is gameobject.Slider {
			// Color
			cursor.add_transform(
				typ: .color,
				easing: easing.linear,
				time: time.Time{last_object.time.end , object.time.start},
				before: last_object.color,
				after: object.color
			)

			// Movement
			mut mover := movers.get_imover() // linear mover

			if (object.time.start - last_object.time.end) >= 50.0 {
				// Use halfcircle for far objects
				mover = &movers.HalfCircleMover{} // Uncomment to use 
			}

			mover.init(mut last_object, mut object, direction)
			direction *= -1 // Invert direction

			for i := mover.time.start; i < mover.time.end; i += offset {
				position := mover.get_point_at(i)
				cursor.add_transform(
					typ: .move, 
					easing: easing.quad_out, 
					time: time.Time{i, i + offset}, 
					before: [last_position.x, last_position.y], 
					after: [position.x, position.y]
				)
				last_position = position
			}

			// Slider movement
			if mut object is gameobject.Slider {
				// Normal movement
				for temp_time := int(object.time.start); temp_time <= int(object.time.end) + offset; temp_time += int(offset) {
					times := int(((temp_time - object.time.start) / object.duration) + 1)
					t_time := (f64(temp_time) - object.time.start - (times - 1) * object.duration)
					rt := object.pixel_length / object.curve.length

					mut pos := vector.Vector2{}
					if (times % 2) == 1 {
						pos = object.curve.point_at(rt * t_time / object.duration)
						last_position = object.curve.point_at(rt * (t_time - offset) / object.duration)
					} else {
						pos = object.curve.point_at((1.0 - t_time / object.duration) * rt)
						last_position = object.curve.point_at((1.0 - (t_time - offset) / object.duration) * rt)
					}
					cursor.add_transform(typ: .move, easing: easing.quad_out, time: time.Time{temp_time, temp_time + offset}, before: [last_position.x, last_position.y], after: [pos.x, pos.y])
				}

				// Dance Movement
				// mut slider_mover := &movers.HalfCircleMover{}
				// slider_mover.init(object.hitcircle, object, direction)
				// slider_mover.time.start = object.time.start
				// slider_mover.time.end = object.time.end
				// slider_mover.start = object.hitcircle.position
				// slider_mover.end = object.end_position
				// slider_mover.middle.x = (slider_mover.start.x + slider_mover.end.x) / 2.0
				// slider_mover.middle.y = (slider_mover.start.y + slider_mover.end.y) / 2.0
				// slider_mover.radius = slider_mover.middle.distance(slider_mover.start)
				// slider_mover.ang = math.atan2(slider_mover.start.y - slider_mover.middle.y, slider_mover.start.x - slider_mover.middle.x)

				// for i := slider_mover.time.start; i < slider_mover.time.end; i += offset {
				// 	position := slider_mover.get_point_at(i)
				// 	cursor.add_transform(
				// 		typ: .move, 
				// 		easing: easing.quad_out, 
				// 		time: time.Time{i, i + offset}, 
				// 		before: [last_position.x, last_position.y], 
				// 		after: [position.x, position.y]
				// 	)
				// 	last_position = position
				// }
			}
		} else if mut object is gameobject.Spinner {
			// oh man here we go agane

			speed := 0.85
			radius := 100.0
			timeframe := 16.6667
			mut rotation := 0.0

			last_position = vector.Vector2{
				math.cos(rotation) * radius + 512.0 / 2.0,
				math.sin(rotation) * radius + 384.0 / 2.0
			}

			for i := object.time.start; i < object.time.end; i += timeframe {
				position := vector.Vector2{
					math.cos(rotation) * radius + 512.0 / 2.0,
					math.sin(rotation) * radius + 384.0 / 2.0
				}

				cursor.add_transform(
					typ: .move, 
					easing: easing.linear, 
					time: time.Time{i, i + timeframe},
					before: [last_position.x, last_position.y],
					after: [position.x, position.y],

				)
				
				rotation += speed
				last_position = position
			}
		}


		last_object = unsafe { object }
	}

	cursor.reset_attributes_based_on_transforms()
}