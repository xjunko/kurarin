module object