module player

pub struct Player {
pub mut:
	name string
}
