module player

pub struct Player {
pub mut:
	player_name string
}
