module graphic

pub const (
	bruh_vertices = [
		f32(288.376), 280.0, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 287.55923, 287.7709, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 287.55923, 287.7709, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 285.14468, 295.20218, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 285.14468, 295.20218, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 281.23782, 301.96906, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 281.23782, 301.96906, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 276.00943, 307.7758, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 276.00943, 307.7758, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 269.688, 312.36856, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 269.688, 312.36856, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 262.5498, 315.5467, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 262.5498, 315.5467, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 254.90686, 317.17126, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 254.90686, 317.17126, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 247.09314, 317.17126, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 247.09314, 317.17126, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 239.45018, 315.5467, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 239.45018, 315.5467, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 232.312, 312.36856, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 232.312, 312.36856, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 225.99057, 307.7758, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 225.99057, 307.7758, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 220.76218, 301.96906, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 220.76218, 301.96906, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 216.85533, 295.20218, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 216.85533, 295.20218, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 214.44075, 287.7709, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 214.44075, 287.7709, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 213.624, 280.0, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 213.624, 280.0, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 214.44075, 272.2291, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 214.44075, 272.2291, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 216.85533, 264.79782, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 216.85533, 264.79782, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 220.76218, 258.03094, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 220.76218, 258.03094, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 225.99057, 252.22421, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 225.99057, 252.22421, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 232.312, 247.63144, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 232.312, 247.63144, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 239.45018, 244.45331, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 239.45018, 244.45331, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 247.09314, 242.82875, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 247.09314, 242.82875, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 254.90686, 242.82875, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 254.90686, 242.82875, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 262.5498, 244.45331, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 262.5498, 244.45331, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 269.688, 247.63144, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 269.688, 247.63144, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 276.00943, 252.22421, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 276.00943, 252.22421, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 281.23782, 258.03094, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 281.23782, 258.03094, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 285.14468, 264.79782, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 285.14468, 264.79782, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 287.55923, 272.2291, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 287.55923, 272.2291, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 288.376, 280.0, 1.0, 251.0, 280.0, 0.0, 0.0, 0.0, 251.0, 280.0, 0.0, 251.0, 280.0, 0.0, 1.0, 0.0, 286.3884, 280.22223, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 285.57162, 287.99313, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 285.57162, 287.99313, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 283.15707, 295.4244, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 283.15707, 295.4244, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 279.2502, 302.19128, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 279.2502, 302.19128, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 274.02182, 307.99802, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 274.02182, 307.99802, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 267.70038, 312.5908, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 267.70038, 312.5908, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 260.5622, 315.76892, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 260.5622, 315.76892, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 252.91924, 317.3935, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 252.91924, 317.3935, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 245.10553, 317.3935, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 245.10553, 317.3935, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 237.46257, 315.76892, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 237.46257, 315.76892, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 230.32439, 312.5908, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 230.32439, 312.5908, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 224.00296, 307.99802, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 224.00296, 307.99802, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 218.77457, 302.19128, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 218.77457, 302.19128, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 214.8677, 295.4244, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 214.8677, 295.4244, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 212.45314, 287.99313, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 212.45314, 287.99313, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 211.63638, 280.22223, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 211.63638, 280.22223, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 212.45314, 272.45132, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 212.45314, 272.45132, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 214.8677, 265.02005, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 214.8677, 265.02005, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 218.77457, 258.25317, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 218.77457, 258.25317, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 224.00296, 252.44646, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 224.00296, 252.44646, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 230.32439, 247.85367, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 230.32439, 247.85367, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 237.46257, 244.67554, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 237.46257, 244.67554, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 245.10553, 243.05098, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 245.10553, 243.05098, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 252.91924, 243.05098, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 252.91924, 243.05098, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 260.5622, 244.67554, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 260.5622, 244.67554, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 267.70038, 247.85367, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 267.70038, 247.85367, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 274.02182, 252.44646, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 274.02182, 252.44646, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 279.2502, 258.25317, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 279.2502, 258.25317, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 283.15707, 265.02005, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 283.15707, 265.02005, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 285.57162, 272.45132, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 285.57162, 272.45132, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 286.3884, 280.22223, 1.0, 249.01239, 280.22223, 0.0, 0.0, 0.0, 249.01239, 280.22223, 0.0, 249.01239, 280.22223, 0.0, 1.0, 0.0, 284.4013, 280.44925, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 283.58456, 288.22015, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 283.58456, 288.22015, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 281.16998, 295.65143, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 281.16998, 295.65143, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 277.26312, 302.4183, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 277.26312, 302.4183, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 272.03473, 308.22504, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 272.03473, 308.22504, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 265.71332, 312.8178, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 265.71332, 312.8178, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 258.57513, 315.99594, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 258.57513, 315.99594, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 250.93217, 317.6205, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 250.93217, 317.6205, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 243.11845, 317.6205, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 243.11845, 317.6205, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 235.4755, 315.99594, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 235.4755, 315.99594, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 228.33731, 312.8178, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 228.33731, 312.8178, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 222.01588, 308.22504, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 222.01588, 308.22504, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 216.78749, 302.4183, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 216.78749, 302.4183, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 212.88063, 295.65143, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 212.88063, 295.65143, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 210.46606, 288.22015, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 210.46606, 288.22015, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 209.6493, 280.44925, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 209.6493, 280.44925, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 210.46606, 272.67834, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 210.46606, 272.67834, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 212.88063, 265.24707, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 212.88063, 265.24707, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 216.78749, 258.4802, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 216.78749, 258.4802, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 222.01588, 252.67348, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 222.01588, 252.67348, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 228.33731, 248.08069, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 228.33731, 248.08069, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 235.4755, 244.90256, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 235.4755, 244.90256, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 243.11845, 243.278, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 243.11845, 243.278, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 250.93217, 243.278, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 250.93217, 243.278, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 258.57513, 244.90256, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 258.57513, 244.90256, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 265.71332, 248.08069, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 265.71332, 248.08069, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 272.03473, 252.67348, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 272.03473, 252.67348, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 277.26312, 258.4802, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 277.26312, 258.4802, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 281.16998, 265.24707, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 281.16998, 265.24707, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 283.58456, 272.67834, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 283.58456, 272.67834, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 284.4013, 280.44925, 1.0, 247.02531, 280.44925, 0.0, 0.0, 0.0, 247.02531, 280.44925, 0.0, 247.02531, 280.44925, 0.0, 1.0, 0.0, 282.4148, 280.68106, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 281.59802, 288.45197, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 281.59802, 288.45197, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 279.18347, 295.88324, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 279.18347, 295.88324, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 275.2766, 302.65012, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 275.2766, 302.65012, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 270.04822, 308.45685, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 270.04822, 308.45685, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 263.7268, 313.04962, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 263.7268, 313.04962, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 256.58862, 316.22775, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 256.58862, 316.22775, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 248.94565, 317.8523, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 248.94565, 317.8523, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 241.13194, 317.8523, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 241.13194, 317.8523, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 233.48897, 316.22775, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 233.48897, 316.22775, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 226.35078, 313.04962, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 226.35078, 313.04962, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 220.02937, 308.45685, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 220.02937, 308.45685, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 214.80098, 302.65012, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 214.80098, 302.65012, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 210.89412, 295.88324, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 210.89412, 295.88324, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 208.47955, 288.45197, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 208.47955, 288.45197, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 207.6628, 280.68106, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 207.6628, 280.68106, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 208.47955, 272.91016, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 208.47955, 272.91016, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 210.89412, 265.47888, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 210.89412, 265.47888, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 214.80098, 258.712, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 214.80098, 258.712, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 220.02937, 252.90527, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 220.02937, 252.90527, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 226.35078, 248.3125, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 226.35078, 248.3125, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 233.48897, 245.13437, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 233.48897, 245.13437, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 241.13194, 243.50981, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 241.13194, 243.50981, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 248.94565, 243.50981, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 248.94565, 243.50981, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 256.58862, 245.13437, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 256.58862, 245.13437, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 263.7268, 248.3125, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 263.7268, 248.3125, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 270.04822, 252.90527, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 270.04822, 252.90527, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 275.2766, 258.712, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 275.2766, 258.712, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 279.18347, 265.47888, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 279.18347, 265.47888, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 281.59802, 272.91016, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 281.59802, 272.91016, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 282.4148, 280.68106, 1.0, 245.03879, 280.68106, 0.0, 0.0, 0.0, 245.03879, 280.68106, 0.0, 245.03879, 280.68106, 0.0, 1.0, 0.0, 280.42883, 280.91766, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 279.6121, 288.68857, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 279.6121, 288.68857, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 277.1975, 296.11984, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 277.1975, 296.11984, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 273.29065, 302.88672, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 273.29065, 302.88672, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 268.06226, 308.69342, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 268.06226, 308.69342, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 261.74084, 313.28622, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 261.74084, 313.28622, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 254.60266, 316.46436, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 254.60266, 316.46436, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 246.95969, 318.0889, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 246.95969, 318.0889, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 239.14598, 318.0889, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 239.14598, 318.0889, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 231.50302, 316.46436, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 231.50302, 316.46436, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 224.36484, 313.28622, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 224.36484, 313.28622, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 218.04341, 308.69342, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 218.04341, 308.69342, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 212.81502, 302.88672, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 212.81502, 302.88672, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 208.90816, 296.11984, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 208.90816, 296.11984, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 206.49359, 288.68857, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 206.49359, 288.68857, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 205.67683, 280.91766, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 205.67683, 280.91766, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 206.49359, 273.14676, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 206.49359, 273.14676, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 208.90816, 265.71545, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 208.90816, 265.71545, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 212.81502, 258.94858, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 212.81502, 258.94858, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 218.04341, 253.14188, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 218.04341, 253.14188, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 224.36484, 248.54909, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 224.36484, 248.54909, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 231.50302, 245.37097, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 231.50302, 245.37097, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 239.14598, 243.7464, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 239.14598, 243.7464, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 246.95969, 243.7464, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 246.95969, 243.7464, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 254.60266, 245.37097, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 254.60266, 245.37097, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 261.74084, 248.54909, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 261.74084, 248.54909, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 268.06226, 253.14188, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 268.06226, 253.14188, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 273.29065, 258.94858, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 273.29065, 258.94858, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 277.1975, 265.71545, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 277.1975, 265.71545, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 279.6121, 273.14676, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 279.6121, 273.14676, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 280.42883, 280.91766, 1.0, 243.05284, 280.91766, 0.0, 0.0, 0.0, 243.05284, 280.91766, 0.0, 243.05284, 280.91766, 0.0, 1.0, 0.0, 278.44345, 281.15903, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 277.6267, 288.92993, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 277.6267, 288.92993, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 275.21213, 296.36124, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 275.21213, 296.36124, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 271.30527, 303.12808, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 271.30527, 303.12808, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 266.07687, 308.9348, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 266.07687, 308.9348, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 259.75546, 313.5276, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 259.75546, 313.5276, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 252.61728, 316.70572, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 252.61728, 316.70572, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 244.97432, 318.3303, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 244.97432, 318.3303, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 237.1606, 318.3303, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 237.1606, 318.3303, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 229.51764, 316.70572, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 229.51764, 316.70572, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 222.37946, 313.5276, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 222.37946, 313.5276, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 216.05803, 308.9348, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 216.05803, 308.9348, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 210.82964, 303.12808, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 210.82964, 303.12808, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 206.92278, 296.36124, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 206.92278, 296.36124, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 204.50821, 288.92993, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 204.50821, 288.92993, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 203.69145, 281.15903, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 203.69145, 281.15903, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 204.50821, 273.38812, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 204.50821, 273.38812, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 206.92278, 265.95685, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 206.92278, 265.95685, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 210.82964, 259.18997, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 210.82964, 259.18997, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 216.05803, 253.38326, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 216.05803, 253.38326, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 222.37946, 248.79047, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 222.37946, 248.79047, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 229.51764, 245.61235, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 229.51764, 245.61235, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 237.1606, 243.9878, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 237.1606, 243.9878, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 244.97432, 243.9878, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 244.97432, 243.9878, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 252.61728, 245.61235, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 252.61728, 245.61235, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 259.75546, 248.79047, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 259.75546, 248.79047, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 266.07687, 253.38326, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 266.07687, 253.38326, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 271.30527, 259.18997, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 271.30527, 259.18997, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 275.21213, 265.95685, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 275.21213, 265.95685, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 277.6267, 273.38812, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 277.6267, 273.38812, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 278.44345, 281.15903, 1.0, 241.06746, 281.15903, 0.0, 0.0, 0.0, 241.06746, 281.15903, 0.0, 241.06746, 281.15903, 0.0, 1.0, 0.0, 276.45865, 281.4052, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 275.6419, 289.17612, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 275.6419, 289.17612, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 273.22733, 296.6074, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 273.22733, 296.6074, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 269.3205, 303.37427, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 269.3205, 303.37427, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 264.0921, 309.18097, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 264.0921, 309.18097, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 257.77066, 313.77377, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 257.77066, 313.77377, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 250.63248, 316.9519, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 250.63248, 316.9519, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 242.98952, 318.57645, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 242.98952, 318.57645, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 235.17581, 318.57645, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 235.17581, 318.57645, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 227.53285, 316.9519, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 227.53285, 316.9519, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 220.39467, 313.77377, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 220.39467, 313.77377, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 214.07324, 309.18097, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 214.07324, 309.18097, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 208.84485, 303.37427, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 208.84485, 303.37427, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 204.93799, 296.6074, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 204.93799, 296.6074, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 202.52342, 289.17612, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 202.52342, 289.17612, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 201.70667, 281.4052, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 201.70667, 281.4052, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 202.52342, 273.6343, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 202.52342, 273.6343, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 204.93799, 266.203, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 204.93799, 266.203, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 208.84485, 259.43613, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 208.84485, 259.43613, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 214.07324, 253.62943, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 214.07324, 253.62943, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 220.39467, 249.03664, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 220.39467, 249.03664, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 227.53285, 245.8585, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 227.53285, 245.8585, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 235.17581, 244.23395, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 235.17581, 244.23395, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 242.98952, 244.23395, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 242.98952, 244.23395, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 250.63248, 245.8585, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 250.63248, 245.8585, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 257.77066, 249.03664, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 257.77066, 249.03664, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 264.0921, 253.62943, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 264.0921, 253.62943, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 269.3205, 259.43613, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 269.3205, 259.43613, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 273.22733, 266.203, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 273.22733, 266.203, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 275.6419, 273.6343, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 275.6419, 273.6343, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 276.45865, 281.4052, 1.0, 239.08266, 281.4052, 0.0, 0.0, 0.0, 239.08266, 281.4052, 0.0, 239.08266, 281.4052, 0.0, 1.0, 0.0, 274.47446, 281.65616, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 273.6577, 289.42706, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 273.6577, 289.42706, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 271.24313, 296.85834, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 271.24313, 296.85834, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 267.3363, 303.6252, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 267.3363, 303.6252, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 262.1079, 309.43192, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 262.1079, 309.43192, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 255.78647, 314.02472, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 255.78647, 314.02472, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 248.64828, 317.20285, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 248.64828, 317.20285, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 241.00533, 318.8274, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 241.00533, 318.8274, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 233.19162, 318.8274, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 233.19162, 318.8274, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 225.54865, 317.20285, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 225.54865, 317.20285, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 218.41048, 314.02472, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 218.41048, 314.02472, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 212.08905, 309.43192, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 212.08905, 309.43192, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 206.86066, 303.6252, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 206.86066, 303.6252, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 202.9538, 296.85834, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 202.9538, 296.85834, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 200.53923, 289.42706, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 200.53923, 289.42706, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 199.72247, 281.65616, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 199.72247, 281.65616, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 200.53923, 273.88525, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 200.53923, 273.88525, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 202.9538, 266.45395, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 202.9538, 266.45395, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 206.86066, 259.68707, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 206.86066, 259.68707, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 212.08905, 253.88037, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 212.08905, 253.88037, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 218.41048, 249.28758, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 218.41048, 249.28758, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 225.54865, 246.10947, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 225.54865, 246.10947, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 233.19162, 244.4849, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 233.19162, 244.4849, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 241.00533, 244.4849, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 241.00533, 244.4849, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 248.64828, 246.10947, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 248.64828, 246.10947, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 255.78647, 249.28758, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 255.78647, 249.28758, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 262.1079, 253.88037, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 262.1079, 253.88037, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 267.3363, 259.68707, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 267.3363, 259.68707, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 271.24313, 266.45395, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 271.24313, 266.45395, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 273.6577, 273.88525, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 273.6577, 273.88525, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 274.47446, 281.65616, 1.0, 237.09846, 281.65616, 0.0, 0.0, 0.0, 237.09846, 281.65616, 0.0, 237.09846, 281.65616, 0.0, 1.0, 0.0, 272.49088, 281.91187, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 271.67413, 289.6828, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 271.67413, 289.6828, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 269.25955, 297.11407, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 269.25955, 297.11407, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 265.35272, 303.88095, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 265.35272, 303.88095, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 260.12433, 309.68765, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 260.12433, 309.68765, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 253.80289, 314.28046, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 253.80289, 314.28046, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 246.6647, 317.45856, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 246.6647, 317.45856, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 239.02174, 319.08313, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 239.02174, 319.08313, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 231.20804, 319.08313, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 231.20804, 319.08313, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 223.56506, 317.45856, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 223.56506, 317.45856, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 216.4269, 314.28046, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 216.4269, 314.28046, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 210.10547, 309.68765, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 210.10547, 309.68765, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 204.87708, 303.88095, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 204.87708, 303.88095, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 200.97021, 297.11407, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 200.97021, 297.11407, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 198.55565, 289.6828, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 198.55565, 289.6828, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 197.73889, 281.91187, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 197.73889, 281.91187, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 198.55565, 274.14096, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 198.55565, 274.14096, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 200.97021, 266.7097, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 200.97021, 266.7097, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 204.87708, 259.9428, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 204.87708, 259.9428, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 210.10547, 254.1361, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 210.10547, 254.1361, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 216.4269, 249.54332, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 216.4269, 249.54332, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 223.56506, 246.36519, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 223.56506, 246.36519, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 231.20804, 244.74063, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 231.20804, 244.74063, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 239.02174, 244.74063, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 239.02174, 244.74063, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 246.6647, 246.36519, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 246.6647, 246.36519, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 253.80289, 249.54332, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 253.80289, 249.54332, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 260.12433, 254.1361, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 260.12433, 254.1361, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 265.35272, 259.9428, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 265.35272, 259.9428, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 269.25955, 266.7097, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 269.25955, 266.7097, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 271.67413, 274.14096, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 271.67413, 274.14096, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 272.49088, 281.91187, 1.0, 235.11488, 281.91187, 0.0, 0.0, 0.0, 235.11488, 281.91187, 0.0, 235.11488, 281.91187, 0.0, 1.0, 0.0, 270.50793, 282.1724, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 269.69116, 289.9433, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 269.69116, 289.9433, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 267.2766, 297.37457, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 267.2766, 297.37457, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 263.36975, 304.14145, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 263.36975, 304.14145, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 258.14136, 309.94818, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 258.14136, 309.94818, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 251.81993, 314.54095, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 251.81993, 314.54095, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 244.68175, 317.7191, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 244.68175, 317.7191, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 237.03879, 319.34363, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 237.03879, 319.34363, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 229.22507, 319.34363, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 229.22507, 319.34363, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 221.5821, 317.7191, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 221.5821, 317.7191, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 214.44392, 314.54095, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 214.44392, 314.54095, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 208.1225, 309.94818, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 208.1225, 309.94818, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 202.8941, 304.14145, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 202.8941, 304.14145, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 198.98726, 297.37457, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 198.98726, 297.37457, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 196.57268, 289.9433, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 196.57268, 289.9433, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 195.75592, 282.1724, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 195.75592, 282.1724, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 196.57268, 274.4015, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 196.57268, 274.4015, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 198.98726, 266.9702, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 198.98726, 266.9702, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 202.8941, 260.20334, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 202.8941, 260.20334, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 208.1225, 254.3966, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 208.1225, 254.3966, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 214.44392, 249.80382, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 214.44392, 249.80382, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 221.5821, 246.6257, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 221.5821, 246.6257, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 229.22507, 245.00114, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 229.22507, 245.00114, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 237.03879, 245.00114, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 237.03879, 245.00114, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 244.68175, 246.6257, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 244.68175, 246.6257, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 251.81993, 249.80382, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 251.81993, 249.80382, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 258.14136, 254.3966, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 258.14136, 254.3966, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 263.36975, 260.20334, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 263.36975, 260.20334, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 267.2766, 266.9702, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 267.2766, 266.9702, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 269.69116, 274.4015, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 269.69116, 274.4015, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 270.50793, 282.1724, 1.0, 233.13193, 282.1724, 0.0, 0.0, 0.0, 233.13193, 282.1724, 0.0, 233.13193, 282.1724, 0.0, 1.0, 0.0, 268.5256, 282.43768, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 267.70883, 290.2086, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 267.70883, 290.2086, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 265.29428, 297.63986, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 265.29428, 297.63986, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 261.38742, 304.40674, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 261.38742, 304.40674, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 256.15903, 310.21347, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 256.15903, 310.21347, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 249.8376, 314.80624, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 249.8376, 314.80624, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 242.69942, 317.98438, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 242.69942, 317.98438, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 235.05646, 319.60892, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 235.05646, 319.60892, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 227.24274, 319.60892, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 227.24274, 319.60892, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 219.59978, 317.98438, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 219.59978, 317.98438, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 212.4616, 314.80624, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 212.4616, 314.80624, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 206.14017, 310.21347, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 206.14017, 310.21347, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 200.91177, 304.40674, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 200.91177, 304.40674, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 197.00493, 297.63986, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 197.00493, 297.63986, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 194.59036, 290.2086, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 194.59036, 290.2086, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 193.7736, 282.43768, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 193.7736, 282.43768, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 194.59036, 274.66678, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 194.59036, 274.66678, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 197.00493, 267.23547, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 197.00493, 267.23547, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 200.91177, 260.46863, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 200.91177, 260.46863, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 206.14017, 254.6619, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 206.14017, 254.6619, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 212.4616, 250.0691, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 212.4616, 250.0691, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 219.59978, 246.89099, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 219.59978, 246.89099, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 227.24274, 245.26642, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 227.24274, 245.26642, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 235.05646, 245.26642, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 235.05646, 245.26642, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 242.69942, 246.89099, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 242.69942, 246.89099, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 249.8376, 250.0691, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 249.8376, 250.0691, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 256.15903, 254.6619, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 256.15903, 254.6619, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 261.38742, 260.46863, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 261.38742, 260.46863, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 265.29428, 267.23547, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 265.29428, 267.23547, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 267.70883, 274.66678, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 267.70883, 274.66678, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 268.5256, 282.43768, 1.0, 231.1496, 282.43768, 0.0, 0.0, 0.0, 231.1496, 282.43768, 0.0, 231.1496, 282.43768, 0.0, 1.0, 0.0, 266.5439, 282.70773, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 265.72717, 290.47864, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 265.72717, 290.47864, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 263.3126, 297.90994, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 263.3126, 297.90994, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 259.40573, 304.6768, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 259.40573, 304.6768, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 254.17734, 310.48352, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 254.17734, 310.48352, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 247.85591, 315.0763, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 247.85591, 315.0763, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 240.71774, 318.25443, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 240.71774, 318.25443, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 233.07477, 319.879, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 233.07477, 319.879, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 225.26106, 319.879, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 225.26106, 319.879, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 217.6181, 318.25443, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 217.6181, 318.25443, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 210.47992, 315.0763, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 210.47992, 315.0763, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 204.1585, 310.48352, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 204.1585, 310.48352, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 198.9301, 304.6768, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 198.9301, 304.6768, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 195.02324, 297.90994, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 195.02324, 297.90994, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 192.60867, 290.47864, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 192.60867, 290.47864, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 191.79192, 282.70773, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 191.79192, 282.70773, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 192.60867, 274.93683, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 192.60867, 274.93683, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 195.02324, 267.50555, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 195.02324, 267.50555, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 198.9301, 260.73868, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 198.9301, 260.73868, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 204.1585, 254.93196, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 204.1585, 254.93196, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 210.47992, 250.33917, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 210.47992, 250.33917, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 217.6181, 247.16106, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 217.6181, 247.16106, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 225.26106, 245.53648, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 225.26106, 245.53648, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 233.07477, 245.53648, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 233.07477, 245.53648, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 240.71774, 247.16106, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 240.71774, 247.16106, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 247.85591, 250.33917, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 247.85591, 250.33917, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 254.17734, 254.93196, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 254.17734, 254.93196, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 259.40573, 260.73868, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 259.40573, 260.73868, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 263.3126, 267.50555, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 263.3126, 267.50555, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 265.72717, 274.93683, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 265.72717, 274.93683, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 266.5439, 282.70773, 1.0, 229.16792, 282.70773, 0.0, 0.0, 0.0, 229.16792, 282.70773, 0.0, 229.16792, 282.70773, 0.0, 1.0, 0.0, 264.5629, 282.98257, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 263.74612, 290.75348, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 263.74612, 290.75348, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 261.33157, 298.18478, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 261.33157, 298.18478, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 257.4247, 304.95163, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 257.4247, 304.95163, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 252.19632, 310.75836, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 252.19632, 310.75836, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 245.8749, 315.35114, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 245.8749, 315.35114, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 238.73671, 318.52927, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 238.73671, 318.52927, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 231.09375, 320.15384, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 231.09375, 320.15384, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 223.28004, 320.15384, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 223.28004, 320.15384, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 215.63707, 318.52927, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 215.63707, 318.52927, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 208.49889, 315.35114, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 208.49889, 315.35114, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 202.17747, 310.75836, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 202.17747, 310.75836, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 196.94908, 304.95163, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 196.94908, 304.95163, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 193.04222, 298.18478, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 193.04222, 298.18478, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 190.62766, 290.75348, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 190.62766, 290.75348, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 189.8109, 282.98257, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 189.8109, 282.98257, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 190.62766, 275.21167, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 190.62766, 275.21167, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 193.04222, 267.7804, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 193.04222, 267.7804, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 196.94908, 261.01352, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 196.94908, 261.01352, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 202.17747, 255.2068, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 202.17747, 255.2068, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 208.49889, 250.61401, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 208.49889, 250.61401, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 215.63707, 247.4359, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 215.63707, 247.4359, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 223.28004, 245.81133, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 223.28004, 245.81133, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 231.09375, 245.81133, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 231.09375, 245.81133, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 238.73671, 247.4359, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 238.73671, 247.4359, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 245.8749, 250.61401, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 245.8749, 250.61401, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 252.19632, 255.2068, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 252.19632, 255.2068, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 257.4247, 261.01352, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 257.4247, 261.01352, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 261.33157, 267.7804, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 261.33157, 267.7804, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 263.74612, 275.21167, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 263.74612, 275.21167, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 264.5629, 282.98257, 1.0, 227.18689, 282.98257, 0.0, 0.0, 0.0, 227.18689, 282.98257, 0.0, 227.18689, 282.98257, 0.0, 1.0, 0.0, 262.58255, 283.2622, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 261.76578, 291.0331, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 261.76578, 291.0331, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 259.3512, 298.4644, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 259.3512, 298.4644, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 255.44435, 305.23126, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 255.44435, 305.23126, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 250.21596, 311.03796, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 250.21596, 311.03796, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 243.89453, 315.63077, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 243.89453, 315.63077, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 236.75635, 318.80887, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 236.75635, 318.80887, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 229.11339, 320.43344, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 229.11339, 320.43344, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 221.29968, 320.43344, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 221.29968, 320.43344, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 213.65672, 318.80887, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 213.65672, 318.80887, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 206.51854, 315.63077, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 206.51854, 315.63077, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 200.19711, 311.03796, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 200.19711, 311.03796, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 194.96872, 305.23126, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 194.96872, 305.23126, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 191.06186, 298.4644, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 191.06186, 298.4644, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 188.6473, 291.0331, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 188.6473, 291.0331, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 187.83054, 283.2622, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 187.83054, 283.2622, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 188.6473, 275.4913, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 188.6473, 275.4913, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 191.06186, 268.06, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 191.06186, 268.06, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 194.96872, 261.29312, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 194.96872, 261.29312, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 200.19711, 255.48642, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 200.19711, 255.48642, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 206.51854, 250.89363, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 206.51854, 250.89363, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 213.65672, 247.7155, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 213.65672, 247.7155, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 221.29968, 246.09094, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 221.29968, 246.09094, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 229.11339, 246.09094, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 229.11339, 246.09094, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 236.75635, 247.7155, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 236.75635, 247.7155, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 243.89453, 250.89363, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 243.89453, 250.89363, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 250.21596, 255.48642, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 250.21596, 255.48642, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 255.44435, 261.29312, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 255.44435, 261.29312, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 259.3512, 268.06, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 259.3512, 268.06, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 261.76578, 275.4913, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 261.76578, 275.4913, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 262.58255, 283.2622, 1.0, 225.20654, 283.2622, 0.0, 0.0, 0.0, 225.20654, 283.2622, 0.0, 225.20654, 283.2622, 0.0, 1.0, 0.0, 260.60284, 283.54657, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 259.7861, 291.31747, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 259.7861, 291.31747, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 257.37152, 298.74878, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 257.37152, 298.74878, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 253.46468, 305.51566, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 253.46468, 305.51566, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 248.23628, 311.32236, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 248.23628, 311.32236, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 241.91486, 315.91513, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 241.91486, 315.91513, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 234.77667, 319.09326, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 234.77667, 319.09326, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 227.13371, 320.71783, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 227.13371, 320.71783, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 219.32, 320.71783, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 219.32, 320.71783, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 211.67703, 319.09326, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 211.67703, 319.09326, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 204.53886, 315.91513, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 204.53886, 315.91513, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 198.21744, 311.32236, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 198.21744, 311.32236, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 192.98904, 305.51566, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 192.98904, 305.51566, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 189.08218, 298.74878, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 189.08218, 298.74878, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 186.66762, 291.31747, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 186.66762, 291.31747, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 185.85086, 283.54657, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 185.85086, 283.54657, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 186.66762, 275.77567, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 186.66762, 275.77567, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 189.08218, 268.3444, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 189.08218, 268.3444, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 192.98904, 261.5775, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 192.98904, 261.5775, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 198.21744, 255.7708, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 198.21744, 255.7708, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 204.53886, 251.17801, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 204.53886, 251.17801, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 211.67703, 247.9999, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 211.67703, 247.9999, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 219.32, 246.37534, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 219.32, 246.37534, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 227.13371, 246.37534, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 227.13371, 246.37534, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 234.77667, 247.9999, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 234.77667, 247.9999, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 241.91486, 251.17801, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 241.91486, 251.17801, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 248.23628, 255.7708, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 248.23628, 255.7708, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 253.46468, 261.5775, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 253.46468, 261.5775, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 257.37152, 268.3444, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 257.37152, 268.3444, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 259.7861, 275.77567, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 259.7861, 275.77567, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 260.60284, 283.54657, 1.0, 223.22685, 283.54657, 0.0, 0.0, 0.0, 223.22685, 283.54657, 0.0, 223.22685, 283.54657, 0.0, 1.0, 0.0, 258.62387, 283.83572, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 257.80713, 291.60663, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 257.80713, 291.60663, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 255.39255, 299.03793, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 255.39255, 299.03793, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 251.48569, 305.8048, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 251.48569, 305.8048, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 246.2573, 311.6115, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 246.2573, 311.6115, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 239.93587, 316.2043, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 239.93587, 316.2043, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 232.79768, 319.38242, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 232.79768, 319.38242, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 225.15472, 321.007, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 225.15472, 321.007, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 217.34102, 321.007, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 217.34102, 321.007, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 209.69806, 319.38242, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 209.69806, 319.38242, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 202.55988, 316.2043, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 202.55988, 316.2043, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 196.23845, 311.6115, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 196.23845, 311.6115, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 191.01006, 305.8048, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 191.01006, 305.8048, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 187.1032, 299.03793, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 187.1032, 299.03793, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 184.68863, 291.60663, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 184.68863, 291.60663, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 183.87187, 283.83572, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 183.87187, 283.83572, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 184.68863, 276.06482, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 184.68863, 276.06482, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 187.1032, 268.63354, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 187.1032, 268.63354, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 191.01006, 261.86667, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 191.01006, 261.86667, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 196.23845, 256.05997, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 196.23845, 256.05997, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 202.55988, 251.46718, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 202.55988, 251.46718, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 209.69806, 248.28905, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 209.69806, 248.28905, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 217.34102, 246.66449, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 217.34102, 246.66449, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 225.15472, 246.66449, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 225.15472, 246.66449, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 232.79768, 248.28905, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 232.79768, 248.28905, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 239.93587, 251.46718, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 239.93587, 251.46718, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 246.2573, 256.05997, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 246.2573, 256.05997, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 251.48569, 261.86667, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 251.48569, 261.86667, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 255.39255, 268.63354, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 255.39255, 268.63354, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 257.80713, 276.06482, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 257.80713, 276.06482, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 258.62387, 283.83572, 1.0, 221.24788, 283.83572, 0.0, 0.0, 0.0, 221.24788, 283.83572, 0.0, 221.24788, 283.83572, 0.0, 1.0, 0.0, 256.6456, 284.12967, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 255.82883, 291.90057, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 255.82883, 291.90057, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 253.41426, 299.33185, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 253.41426, 299.33185, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 249.5074, 306.09872, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 249.5074, 306.09872, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 244.279, 311.90546, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 244.279, 311.90546, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 237.9576, 316.49823, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 237.9576, 316.49823, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 230.81941, 319.67636, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 230.81941, 319.67636, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 223.17644, 321.3009, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 223.17644, 321.3009, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 215.36273, 321.3009, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 215.36273, 321.3009, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 207.71977, 319.67636, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 207.71977, 319.67636, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 200.58159, 316.49823, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 200.58159, 316.49823, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 194.26016, 311.90546, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 194.26016, 311.90546, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 189.03177, 306.09872, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 189.03177, 306.09872, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 185.12491, 299.33185, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 185.12491, 299.33185, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 182.71034, 291.90057, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 182.71034, 291.90057, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 181.89359, 284.12967, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 181.89359, 284.12967, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 182.71034, 276.35876, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 182.71034, 276.35876, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 185.12491, 268.92746, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 185.12491, 268.92746, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 189.03177, 262.1606, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 189.03177, 262.1606, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 194.26016, 256.35388, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 194.26016, 256.35388, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 200.58159, 251.7611, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 200.58159, 251.7611, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 207.71977, 248.58298, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 207.71977, 248.58298, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 215.36273, 246.9584, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 215.36273, 246.9584, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 223.17644, 246.9584, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 223.17644, 246.9584, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 230.81941, 248.58298, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 230.81941, 248.58298, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 237.9576, 251.7611, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 237.9576, 251.7611, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 244.279, 256.35388, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 244.279, 256.35388, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 249.5074, 262.1606, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 249.5074, 262.1606, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 253.41426, 268.92746, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 253.41426, 268.92746, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 255.82883, 276.35876, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 255.82883, 276.35876, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 256.6456, 284.12967, 1.0, 219.26959, 284.12967, 0.0, 0.0, 0.0, 219.26959, 284.12967, 0.0, 219.26959, 284.12967, 0.0, 1.0, 0.0, 254.66801, 284.42834, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 253.85126, 292.19925, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 253.85126, 292.19925, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 251.43669, 299.63055, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 251.43669, 299.63055, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 247.52983, 306.3974, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 247.52983, 306.3974, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 242.30144, 312.20413, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 242.30144, 312.20413, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 235.98003, 316.7969, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 235.98003, 316.7969, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 228.84184, 319.97504, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 228.84184, 319.97504, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 221.19887, 321.5996, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 221.19887, 321.5996, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 213.38516, 321.5996, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 213.38516, 321.5996, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 205.7422, 319.97504, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 205.7422, 319.97504, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 198.60402, 316.7969, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 198.60402, 316.7969, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 192.2826, 312.20413, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 192.2826, 312.20413, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 187.0542, 306.3974, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 187.0542, 306.3974, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 183.14734, 299.63055, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 183.14734, 299.63055, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 180.73277, 292.19925, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 180.73277, 292.19925, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 179.91602, 284.42834, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 179.91602, 284.42834, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 180.73277, 276.65744, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 180.73277, 276.65744, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 183.14734, 269.22617, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 183.14734, 269.22617, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 187.0542, 262.4593, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 187.0542, 262.4593, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 192.2826, 256.65256, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 192.2826, 256.65256, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 198.60402, 252.05978, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 198.60402, 252.05978, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 205.7422, 248.88167, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 205.7422, 248.88167, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 213.38516, 247.2571, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 213.38516, 247.2571, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 221.19887, 247.2571, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 221.19887, 247.2571, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 228.84184, 248.88167, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 228.84184, 248.88167, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 235.98003, 252.05978, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 235.98003, 252.05978, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 242.30144, 256.65256, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 242.30144, 256.65256, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 247.52983, 262.4593, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 247.52983, 262.4593, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 251.43669, 269.22617, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 251.43669, 269.22617, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 253.85126, 276.65744, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 253.85126, 276.65744, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 254.66801, 284.42834, 1.0, 217.29202, 284.42834, 0.0, 0.0, 0.0, 217.29202, 284.42834, 0.0, 217.29202, 284.42834, 0.0, 1.0, 0.0, 252.69118, 284.7318, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 251.87442, 292.50272, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 251.87442, 292.50272, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 249.45985, 299.934, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 249.45985, 299.934, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 245.553, 306.70087, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 245.553, 306.70087, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 240.3246, 312.5076, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 240.3246, 312.5076, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 234.00317, 317.10037, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 234.00317, 317.10037, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 226.86499, 320.2785, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 226.86499, 320.2785, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 219.22203, 321.90305, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 219.22203, 321.90305, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 211.40833, 321.90305, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 211.40833, 321.90305, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 203.76535, 320.2785, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 203.76535, 320.2785, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 196.62718, 317.10037, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 196.62718, 317.10037, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 190.30576, 312.5076, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 190.30576, 312.5076, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 185.07736, 306.70087, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 185.07736, 306.70087, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 181.1705, 299.934, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 181.1705, 299.934, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 178.75594, 292.50272, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 178.75594, 292.50272, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 177.93918, 284.7318, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 177.93918, 284.7318, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 178.75594, 276.9609, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 178.75594, 276.9609, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 181.1705, 269.52963, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 181.1705, 269.52963, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 185.07736, 262.76276, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 185.07736, 262.76276, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 190.30576, 256.95602, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 190.30576, 256.95602, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 196.62718, 252.36325, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 196.62718, 252.36325, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 203.76535, 249.18512, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 203.76535, 249.18512, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 211.40833, 247.56056, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 211.40833, 247.56056, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 219.22203, 247.56056, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 219.22203, 247.56056, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 226.86499, 249.18512, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 226.86499, 249.18512, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 234.00317, 252.36325, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 234.00317, 252.36325, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 240.3246, 256.95602, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 240.3246, 256.95602, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 245.553, 262.76276, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 245.553, 262.76276, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 249.45985, 269.52963, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 249.45985, 269.52963, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 251.87442, 276.9609, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 251.87442, 276.9609, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 252.69118, 284.7318, 1.0, 215.31517, 284.7318, 0.0, 0.0, 0.0, 215.31517, 284.7318, 0.0, 215.31517, 284.7318, 0.0, 1.0, 0.0, 250.71507, 285.04004, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 249.89832, 292.81094, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 249.89832, 292.81094, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 247.48375, 300.24222, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 247.48375, 300.24222, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 243.57689, 307.0091, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 243.57689, 307.0091, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 238.3485, 312.8158, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 238.3485, 312.8158, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 232.02707, 317.4086, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 232.02707, 317.4086, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 224.88889, 320.58673, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 224.88889, 320.58673, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 217.24593, 322.21127, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 217.24593, 322.21127, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 209.4322, 322.21127, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 209.4322, 322.21127, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 201.78925, 320.58673, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 201.78925, 320.58673, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 194.65106, 317.4086, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 194.65106, 317.4086, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 188.32964, 312.8158, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 188.32964, 312.8158, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 183.10124, 307.0091, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 183.10124, 307.0091, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 179.1944, 300.24222, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 179.1944, 300.24222, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 176.77983, 292.81094, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 176.77983, 292.81094, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 175.96307, 285.04004, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 175.96307, 285.04004, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 176.77983, 277.26913, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 176.77983, 277.26913, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 179.1944, 269.83783, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 179.1944, 269.83783, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 183.10124, 263.07095, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 183.10124, 263.07095, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 188.32964, 257.26425, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 188.32964, 257.26425, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 194.65106, 252.67146, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 194.65106, 252.67146, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 201.78925, 249.49335, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 201.78925, 249.49335, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 209.4322, 247.86877, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 209.4322, 247.86877, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 217.24593, 247.86877, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 217.24593, 247.86877, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 224.88889, 249.49335, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 224.88889, 249.49335, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 232.02707, 252.67146, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 232.02707, 252.67146, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 238.3485, 257.26425, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 238.3485, 257.26425, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 243.57689, 263.07095, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 243.57689, 263.07095, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 247.48375, 269.83783, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 247.48375, 269.83783, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 249.89832, 277.26913, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 249.89832, 277.26913, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 250.71507, 285.04004, 1.0, 213.33907, 285.04004, 0.0, 0.0, 0.0, 213.33907, 285.04004, 0.0, 213.33907, 285.04004, 0.0, 1.0, 0.0, 248.73972, 285.35303, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 247.92296, 293.12393, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 247.92296, 293.12393, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 245.50839, 300.5552, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 245.50839, 300.5552, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 241.60153, 307.32208, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 241.60153, 307.32208, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 236.37314, 313.12878, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 236.37314, 313.12878, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 230.05171, 317.7216, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 230.05171, 317.7216, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 222.91353, 320.8997, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 222.91353, 320.8997, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 215.27057, 322.52426, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 215.27057, 322.52426, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 207.45685, 322.52426, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 207.45685, 322.52426, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 199.81389, 320.8997, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 199.81389, 320.8997, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 192.6757, 317.7216, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 192.6757, 317.7216, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 186.35428, 313.12878, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 186.35428, 313.12878, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 181.12589, 307.32208, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 181.12589, 307.32208, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 177.21904, 300.5552, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 177.21904, 300.5552, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 174.80446, 293.12393, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 174.80446, 293.12393, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 173.98772, 285.35303, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 173.98772, 285.35303, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 174.80446, 277.5821, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 174.80446, 277.5821, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 177.21904, 270.15082, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 177.21904, 270.15082, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 181.12589, 263.38394, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 181.12589, 263.38394, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 186.35428, 257.57724, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 186.35428, 257.57724, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 192.6757, 252.98445, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 192.6757, 252.98445, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 199.81389, 249.80632, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 199.81389, 249.80632, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 207.45685, 248.18176, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 207.45685, 248.18176, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 215.27057, 248.18176, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 215.27057, 248.18176, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 222.91353, 249.80632, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 222.91353, 249.80632, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 230.05171, 252.98445, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 230.05171, 252.98445, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 236.37314, 257.57724, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 236.37314, 257.57724, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 241.60153, 263.38394, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 241.60153, 263.38394, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 245.50839, 270.15082, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 245.50839, 270.15082, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 247.92296, 277.5821, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 247.92296, 277.5821, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 248.73972, 285.35303, 1.0, 211.36371, 285.35303, 0.0, 0.0, 0.0, 211.36371, 285.35303, 0.0, 211.36371, 285.35303, 0.0, 1.0, 0.0, 246.7651, 285.67075, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 245.94835, 293.44165, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 245.94835, 293.44165, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 243.53378, 300.87296, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 243.53378, 300.87296, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 239.62694, 307.6398, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 239.62694, 307.6398, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 234.39854, 313.44653, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 234.39854, 313.44653, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 228.07712, 318.0393, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 228.07712, 318.0393, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 220.93893, 321.21744, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 220.93893, 321.21744, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 213.29597, 322.842, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 213.29597, 322.842, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 205.48225, 322.842, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 205.48225, 322.842, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 197.8393, 321.21744, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 197.8393, 321.21744, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 190.70111, 318.0393, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 190.70111, 318.0393, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 184.37968, 313.44653, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 184.37968, 313.44653, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 179.15129, 307.6398, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 179.15129, 307.6398, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 175.24443, 300.87296, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 175.24443, 300.87296, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 172.82986, 293.44165, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 172.82986, 293.44165, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 172.0131, 285.67075, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 172.0131, 285.67075, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 172.82986, 277.89984, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 172.82986, 277.89984, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 175.24443, 270.46857, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 175.24443, 270.46857, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 179.15129, 263.7017, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 179.15129, 263.7017, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 184.37968, 257.89496, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 184.37968, 257.89496, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 190.70111, 253.30219, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 190.70111, 253.30219, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 197.8393, 250.12407, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 197.8393, 250.12407, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 205.48225, 248.4995, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 205.48225, 248.4995, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 213.29597, 248.4995, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 213.29597, 248.4995, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 220.93893, 250.12407, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 220.93893, 250.12407, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 228.07712, 253.30219, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 228.07712, 253.30219, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 234.39854, 257.89496, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 234.39854, 257.89496, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 239.62694, 263.7017, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 239.62694, 263.7017, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 243.53378, 270.46857, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 243.53378, 270.46857, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 245.94835, 277.89984, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 245.94835, 277.89984, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 246.7651, 285.67075, 1.0, 209.38911, 285.67075, 0.0, 0.0, 0.0, 209.38911, 285.67075, 0.0, 209.38911, 285.67075, 0.0, 1.0, 0.0, 244.79129, 285.99326, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 243.97453, 293.76416, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 243.97453, 293.76416, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 241.55997, 301.19543, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 241.55997, 301.19543, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 237.6531, 307.9623, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 237.6531, 307.9623, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 232.42471, 313.76904, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 232.42471, 313.76904, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 226.10329, 318.36182, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 226.10329, 318.36182, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 218.9651, 321.53995, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 218.9651, 321.53995, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 211.32214, 323.1645, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 211.32214, 323.1645, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 203.50842, 323.1645, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 203.50842, 323.1645, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 195.86546, 321.53995, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 195.86546, 321.53995, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 188.72728, 318.36182, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 188.72728, 318.36182, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 182.40585, 313.76904, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 182.40585, 313.76904, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 177.17746, 307.9623, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 177.17746, 307.9623, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 173.27061, 301.19543, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 173.27061, 301.19543, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 170.85603, 293.76416, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 170.85603, 293.76416, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 170.03929, 285.99326, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 170.03929, 285.99326, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 170.85603, 278.22235, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 170.85603, 278.22235, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 173.27061, 270.79108, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 173.27061, 270.79108, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 177.17746, 264.0242, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 177.17746, 264.0242, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 182.40585, 258.21747, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 182.40585, 258.21747, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 188.72728, 253.6247, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 188.72728, 253.6247, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 195.86546, 250.44656, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 195.86546, 250.44656, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 203.50842, 248.822, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 203.50842, 248.822, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 211.32214, 248.822, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 211.32214, 248.822, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 218.9651, 250.44656, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 218.9651, 250.44656, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 226.10329, 253.6247, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 226.10329, 253.6247, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 232.42471, 258.21747, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 232.42471, 258.21747, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 237.6531, 264.0242, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 237.6531, 264.0242, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 241.55997, 270.79108, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 241.55997, 270.79108, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 243.97453, 278.22235, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 243.97453, 278.22235, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 244.79129, 285.99326, 1.0, 207.41528, 285.99326, 0.0, 0.0, 0.0, 207.41528, 285.99326, 0.0, 207.41528, 285.99326, 0.0, 1.0, 0.0, 242.81824, 286.3205, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 242.00148, 294.09143, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 242.00148, 294.09143, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 239.58691, 301.5227, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 239.58691, 301.5227, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 235.68005, 308.28958, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 235.68005, 308.28958, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 230.45166, 314.09628, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 230.45166, 314.09628, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 224.13023, 318.6891, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 224.13023, 318.6891, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 216.99207, 321.8672, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 216.99207, 321.8672, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 209.34909, 323.49176, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 209.34909, 323.49176, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 201.53539, 323.49176, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 201.53539, 323.49176, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 193.89243, 321.8672, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 193.89243, 321.8672, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 186.75424, 318.6891, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 186.75424, 318.6891, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 180.43282, 314.09628, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 180.43282, 314.09628, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 175.20442, 308.28958, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 175.20442, 308.28958, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 171.29756, 301.5227, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 171.29756, 301.5227, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 168.883, 294.09143, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 168.883, 294.09143, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 168.06624, 286.3205, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 168.06624, 286.3205, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 168.883, 278.5496, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 168.883, 278.5496, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 171.29756, 271.11832, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 171.29756, 271.11832, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 175.20442, 264.35144, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 175.20442, 264.35144, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 180.43282, 258.54474, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 180.43282, 258.54474, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 186.75424, 253.95195, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 186.75424, 253.95195, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 193.89243, 250.77382, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 193.89243, 250.77382, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 201.53539, 249.14926, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 201.53539, 249.14926, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 209.34909, 249.14926, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 209.34909, 249.14926, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 216.99207, 250.77382, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 216.99207, 250.77382, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 224.13023, 253.95195, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 224.13023, 253.95195, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 230.45166, 258.54474, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 230.45166, 258.54474, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 235.68005, 264.35144, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 235.68005, 264.35144, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 239.58691, 271.11832, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 239.58691, 271.11832, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 242.00148, 278.5496, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 242.00148, 278.5496, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 242.81824, 286.3205, 1.0, 205.44225, 286.3205, 0.0, 0.0, 0.0, 205.44225, 286.3205, 0.0, 205.44225, 286.3205, 0.0, 1.0, 0.0, 240.846, 286.65253, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 240.02924, 294.42343, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 240.02924, 294.42343, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 237.61467, 301.8547, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 237.61467, 301.8547, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 233.70781, 308.62158, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 233.70781, 308.62158, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 228.47942, 314.4283, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 228.47942, 314.4283, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 222.15799, 319.0211, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 222.15799, 319.0211, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 215.0198, 322.19922, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 215.0198, 322.19922, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 207.37685, 323.82376, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 207.37685, 323.82376, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 199.56314, 323.82376, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 199.56314, 323.82376, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 191.92017, 322.19922, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 191.92017, 322.19922, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 184.782, 319.0211, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 184.782, 319.0211, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 178.46057, 314.4283, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 178.46057, 314.4283, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 173.23218, 308.62158, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 173.23218, 308.62158, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 169.32532, 301.8547, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 169.32532, 301.8547, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 166.91075, 294.42343, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 166.91075, 294.42343, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 166.094, 286.65253, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 166.094, 286.65253, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 166.91075, 278.88162, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 166.91075, 278.88162, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 169.32532, 271.45032, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 169.32532, 271.45032, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 173.23218, 264.68347, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 173.23218, 264.68347, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 178.46057, 258.87674, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 178.46057, 258.87674, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 184.782, 254.28395, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 184.782, 254.28395, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 191.92017, 251.10583, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 191.92017, 251.10583, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 199.56314, 249.48128, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 199.56314, 249.48128, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 207.37685, 249.48128, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 207.37685, 249.48128, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 215.0198, 251.10583, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 215.0198, 251.10583, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 222.15799, 254.28395, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 222.15799, 254.28395, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 228.47942, 258.87674, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 228.47942, 258.87674, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 233.70781, 264.68347, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 233.70781, 264.68347, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 237.61467, 271.45032, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 237.61467, 271.45032, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 240.02924, 278.88162, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 240.02924, 278.88162, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 240.846, 286.65253, 1.0, 203.46999, 286.65253, 0.0, 0.0, 0.0, 203.46999, 286.65253, 0.0, 203.46999, 286.65253, 0.0, 1.0, 0.0, 238.87454, 286.9893, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 238.0578, 294.7602, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 238.0578, 294.7602, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 235.64322, 302.19147, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 235.64322, 302.19147, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 231.73637, 308.95834, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 231.73637, 308.95834, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 226.50798, 314.76508, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 226.50798, 314.76508, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 220.18655, 319.35785, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 220.18655, 319.35785, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 213.04837, 322.53598, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 213.04837, 322.53598, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 205.40541, 324.16052, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 205.40541, 324.16052, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 197.59169, 324.16052, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 197.59169, 324.16052, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 189.94873, 322.53598, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 189.94873, 322.53598, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 182.81055, 319.35785, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 182.81055, 319.35785, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 176.48912, 314.76508, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 176.48912, 314.76508, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 171.26073, 308.95834, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 171.26073, 308.95834, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 167.35387, 302.19147, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 167.35387, 302.19147, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 164.9393, 294.7602, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 164.9393, 294.7602, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 164.12254, 286.9893, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 164.12254, 286.9893, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 164.9393, 279.21838, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 164.9393, 279.21838, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 167.35387, 271.7871, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 167.35387, 271.7871, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 171.26073, 265.02023, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 171.26073, 265.02023, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 176.48912, 259.2135, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 176.48912, 259.2135, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 182.81055, 254.62071, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 182.81055, 254.62071, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 189.94873, 251.4426, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 189.94873, 251.4426, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 197.59169, 249.81804, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 197.59169, 249.81804, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 205.40541, 249.81804, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 205.40541, 249.81804, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 213.04837, 251.4426, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 213.04837, 251.4426, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 220.18655, 254.62071, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 220.18655, 254.62071, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 226.50798, 259.2135, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 226.50798, 259.2135, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 231.73637, 265.02023, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 231.73637, 265.02023, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 235.64322, 271.7871, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 235.64322, 271.7871, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 238.0578, 279.21838, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 238.0578, 279.21838, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 238.87454, 286.9893, 1.0, 201.49855, 286.9893, 0.0, 0.0, 0.0, 201.49855, 286.9893, 0.0, 201.49855, 286.9893, 0.0, 1.0, 0.0, 236.90392, 287.3308, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 236.08717, 295.1017, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 236.08717, 295.1017, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 233.67259, 302.533, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 233.67259, 302.533, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 229.76575, 309.29987, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 229.76575, 309.29987, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 224.53735, 315.10657, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 224.53735, 315.10657, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 218.21593, 319.69937, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 218.21593, 319.69937, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 211.07774, 322.87747, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 211.07774, 322.87747, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 203.43478, 324.50204, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 203.43478, 324.50204, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 195.62106, 324.50204, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 195.62106, 324.50204, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 187.9781, 322.87747, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 187.9781, 322.87747, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 180.83992, 319.69937, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 180.83992, 319.69937, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 174.5185, 315.10657, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 174.5185, 315.10657, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 169.2901, 309.29987, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 169.2901, 309.29987, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 165.38326, 302.533, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 165.38326, 302.533, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 162.96867, 295.1017, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 162.96867, 295.1017, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 162.15192, 287.3308, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 162.15192, 287.3308, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 162.96867, 279.55988, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 162.96867, 279.55988, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 165.38326, 272.1286, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 165.38326, 272.1286, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 169.2901, 265.36172, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 169.2901, 265.36172, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 174.5185, 259.55502, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 174.5185, 259.55502, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 180.83992, 254.96223, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 180.83992, 254.96223, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 187.9781, 251.7841, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 187.9781, 251.7841, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 195.62106, 250.15955, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 195.62106, 250.15955, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 203.43478, 250.15955, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 203.43478, 250.15955, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 211.07774, 251.7841, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 211.07774, 251.7841, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 218.21593, 254.96223, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 218.21593, 254.96223, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 224.53735, 259.55502, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 224.53735, 259.55502, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 229.76575, 265.36172, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 229.76575, 265.36172, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 233.67259, 272.1286, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 233.67259, 272.1286, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 236.08717, 279.55988, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 236.08717, 279.55988, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 236.90392, 287.3308, 1.0, 199.52792, 287.3308, 0.0, 0.0, 0.0, 199.52792, 287.3308, 0.0, 199.52792, 287.3308, 0.0, 1.0, 0.0, 234.93413, 287.67706, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 234.11737, 295.44797, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 234.11737, 295.44797, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 231.7028, 302.87924, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 231.7028, 302.87924, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 227.79594, 309.64612, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 227.79594, 309.64612, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 222.56755, 315.45285, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 222.56755, 315.45285, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 216.24612, 320.04562, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 216.24612, 320.04562, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 209.10794, 323.22375, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 209.10794, 323.22375, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 201.46498, 324.8483, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 201.46498, 324.8483, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 193.65128, 324.8483, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 193.65128, 324.8483, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 186.0083, 323.22375, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 186.0083, 323.22375, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 178.87013, 320.04562, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 178.87013, 320.04562, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 172.5487, 315.45285, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 172.5487, 315.45285, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 167.32031, 309.64612, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 167.32031, 309.64612, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 163.41345, 302.87924, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 163.41345, 302.87924, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 160.99889, 295.44797, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 160.99889, 295.44797, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 160.18213, 287.67706, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 160.18213, 287.67706, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 160.99889, 279.90616, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 160.99889, 279.90616, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 163.41345, 272.47488, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 163.41345, 272.47488, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 167.32031, 265.708, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 167.32031, 265.708, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 172.5487, 259.90128, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 172.5487, 259.90128, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 178.87013, 255.30849, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 178.87013, 255.30849, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 186.0083, 252.13037, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 186.0083, 252.13037, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 193.65128, 250.50581, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 193.65128, 250.50581, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 201.46498, 250.50581, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 201.46498, 250.50581, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 209.10794, 252.13037, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 209.10794, 252.13037, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 216.24612, 255.30849, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 216.24612, 255.30849, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 222.56755, 259.90128, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 222.56755, 259.90128, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 227.79594, 265.708, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 227.79594, 265.708, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 231.7028, 272.47488, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 231.7028, 272.47488, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 234.11737, 279.90616, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 234.11737, 279.90616, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 234.93413, 287.67706, 1.0, 197.55812, 287.67706, 0.0, 0.0, 0.0, 197.55812, 287.67706, 0.0, 197.55812, 287.67706, 0.0, 1.0, 0.0, 232.96516, 288.02808, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 232.1484, 295.79898, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 232.1484, 295.79898, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 229.73384, 303.23026, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 229.73384, 303.23026, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 225.82698, 309.99713, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 225.82698, 309.99713, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 220.59859, 315.80383, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 220.59859, 315.80383, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 214.27718, 320.39664, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 214.27718, 320.39664, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 207.13899, 323.57477, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 207.13899, 323.57477, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 199.49602, 325.1993, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 199.49602, 325.1993, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 191.68231, 325.1993, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 191.68231, 325.1993, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 184.03935, 323.57477, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 184.03935, 323.57477, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 176.90117, 320.39664, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 176.90117, 320.39664, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 170.57974, 315.80383, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 170.57974, 315.80383, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 165.35135, 309.99713, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 165.35135, 309.99713, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 161.44449, 303.23026, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 161.44449, 303.23026, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 159.02992, 295.79898, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 159.02992, 295.79898, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 158.21317, 288.02808, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 158.21317, 288.02808, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 159.02992, 280.25717, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 159.02992, 280.25717, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 161.44449, 272.82587, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 161.44449, 272.82587, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 165.35135, 266.059, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 165.35135, 266.059, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 170.57974, 260.2523, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 170.57974, 260.2523, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 176.90117, 255.6595, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 176.90117, 255.6595, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 184.03935, 252.48138, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 184.03935, 252.48138, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 191.68231, 250.85681, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 191.68231, 250.85681, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 199.49602, 250.85681, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 199.49602, 250.85681, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 207.13899, 252.48138, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 207.13899, 252.48138, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 214.27718, 255.6595, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 214.27718, 255.6595, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 220.59859, 260.2523, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 220.59859, 260.2523, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 225.82698, 266.059, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 225.82698, 266.059, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 229.73384, 272.82587, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 229.73384, 272.82587, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 232.1484, 280.25717, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 232.1484, 280.25717, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 232.96516, 288.02808, 1.0, 195.58917, 288.02808, 0.0, 0.0, 0.0, 195.58917, 288.02808, 0.0, 195.58917, 288.02808, 0.0, 1.0, 0.0, 230.99707, 288.38382, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 230.18031, 296.15472, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 230.18031, 296.15472, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 227.76573, 303.586, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 227.76573, 303.586, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 223.85889, 310.35287, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 223.85889, 310.35287, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 218.6305, 316.1596, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 218.6305, 316.1596, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 212.30907, 320.75238, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 212.30907, 320.75238, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 205.17088, 323.9305, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 205.17088, 323.9305, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 197.52792, 325.55508, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 197.52792, 325.55508, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 189.7142, 325.55508, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 189.7142, 325.55508, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 182.07124, 323.9305, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 182.07124, 323.9305, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 174.93306, 320.75238, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 174.93306, 320.75238, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 168.61163, 316.1596, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 168.61163, 316.1596, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 163.38324, 310.35287, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 163.38324, 310.35287, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 159.4764, 303.586, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 159.4764, 303.586, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 157.06181, 296.15472, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 157.06181, 296.15472, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 156.24506, 288.38382, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 156.24506, 288.38382, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 157.06181, 280.6129, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 157.06181, 280.6129, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 159.4764, 273.18164, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 159.4764, 273.18164, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 163.38324, 266.41476, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 163.38324, 266.41476, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 168.61163, 260.60803, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 168.61163, 260.60803, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 174.93306, 256.01526, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 174.93306, 256.01526, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 182.07124, 252.83713, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 182.07124, 252.83713, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 189.7142, 251.21257, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 189.7142, 251.21257, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 197.52792, 251.21257, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 197.52792, 251.21257, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 205.17088, 252.83713, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 205.17088, 252.83713, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 212.30907, 256.01526, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 212.30907, 256.01526, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 218.6305, 260.60803, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 218.6305, 260.60803, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 223.85889, 266.41476, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 223.85889, 266.41476, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 227.76573, 273.18164, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 227.76573, 273.18164, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 230.18031, 280.6129, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 230.18031, 280.6129, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 230.99707, 288.38382, 1.0, 193.62106, 288.38382, 0.0, 0.0, 0.0, 193.62106, 288.38382, 0.0, 193.62106, 288.38382, 0.0, 1.0, 0.0, 229.02982, 288.74432, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 228.21306, 296.51523, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 228.21306, 296.51523, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 225.7985, 303.9465, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 225.7985, 303.9465, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 221.89165, 310.71338, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 221.89165, 310.71338, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 216.66325, 316.52008, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 216.66325, 316.52008, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 210.34183, 321.11288, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 210.34183, 321.11288, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 203.20364, 324.29102, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 203.20364, 324.29102, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 195.56068, 325.91556, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 195.56068, 325.91556, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 187.74696, 325.91556, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 187.74696, 325.91556, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 180.104, 324.29102, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 180.104, 324.29102, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 172.96582, 321.11288, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 172.96582, 321.11288, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 166.6444, 316.52008, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 166.6444, 316.52008, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 161.416, 310.71338, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 161.416, 310.71338, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 157.50914, 303.9465, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 157.50914, 303.9465, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 155.09457, 296.51523, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 155.09457, 296.51523, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 154.27782, 288.74432, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 154.27782, 288.74432, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 155.09457, 280.97342, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 155.09457, 280.97342, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 157.50914, 273.5421, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 157.50914, 273.5421, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 161.416, 266.77524, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 161.416, 266.77524, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 166.6444, 260.96854, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 166.6444, 260.96854, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 172.96582, 256.37576, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 172.96582, 256.37576, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 180.104, 253.19763, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 180.104, 253.19763, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 187.74696, 251.57306, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 187.74696, 251.57306, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 195.56068, 251.57306, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 195.56068, 251.57306, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 203.20364, 253.19763, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 203.20364, 253.19763, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 210.34183, 256.37576, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 210.34183, 256.37576, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 216.66325, 260.96854, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 216.66325, 260.96854, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 221.89165, 266.77524, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 221.89165, 266.77524, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 225.7985, 273.5421, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 225.7985, 273.5421, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 228.21306, 280.97342, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 228.21306, 280.97342, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 229.02982, 288.74432, 1.0, 191.65382, 288.74432, 0.0, 0.0, 0.0, 191.65382, 288.74432, 0.0, 191.65382, 288.74432, 0.0, 1.0, 0.0, 227.06345, 289.10956, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 226.2467, 296.88046, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 226.2467, 296.88046, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 223.83212, 304.31174, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 223.83212, 304.31174, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 219.92528, 311.0786, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 219.92528, 311.0786, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 214.69688, 316.8853, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 214.69688, 316.8853, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 208.37546, 321.47812, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 208.37546, 321.47812, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 201.23727, 324.65625, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 201.23727, 324.65625, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 193.59431, 326.2808, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 193.59431, 326.2808, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 185.7806, 326.2808, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 185.7806, 326.2808, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 178.13763, 324.65625, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 178.13763, 324.65625, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 170.99945, 321.47812, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 170.99945, 321.47812, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 164.67802, 316.8853, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 164.67802, 316.8853, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 159.44963, 311.0786, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 159.44963, 311.0786, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 155.54279, 304.31174, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 155.54279, 304.31174, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 153.1282, 296.88046, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 153.1282, 296.88046, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 152.31145, 289.10956, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 152.31145, 289.10956, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 153.1282, 281.33865, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 153.1282, 281.33865, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 155.54279, 273.90735, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 155.54279, 273.90735, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 159.44963, 267.14047, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 159.44963, 267.14047, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 164.67802, 261.33377, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 164.67802, 261.33377, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 170.99945, 256.741, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 170.99945, 256.741, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 178.13763, 253.56287, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 178.13763, 253.56287, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 185.7806, 251.9383, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 185.7806, 251.9383, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 193.59431, 251.9383, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 193.59431, 251.9383, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 201.23727, 253.56287, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 201.23727, 253.56287, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 208.37546, 256.741, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 208.37546, 256.741, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 214.69688, 261.33377, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 214.69688, 261.33377, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 219.92528, 267.14047, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 219.92528, 267.14047, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 223.83212, 273.90735, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 223.83212, 273.90735, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 226.2467, 281.33865, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 226.2467, 281.33865, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 227.06345, 289.10956, 1.0, 189.68745, 289.10956, 0.0, 0.0, 0.0, 189.68745, 289.10956, 0.0, 189.68745, 289.10956, 0.0, 1.0, 0.0, 225.09798, 289.47952, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 224.28122, 297.25043, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 224.28122, 297.25043, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 221.86665, 304.6817, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 221.86665, 304.6817, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 217.9598, 311.44858, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 217.9598, 311.44858, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 212.7314, 317.2553, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 212.7314, 317.2553, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 206.40997, 321.84808, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 206.40997, 321.84808, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 199.27179, 325.0262, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 199.27179, 325.0262, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 191.62883, 326.6508, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 191.62883, 326.6508, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 183.81511, 326.6508, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 183.81511, 326.6508, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 176.17215, 325.0262, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 176.17215, 325.0262, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 169.03397, 321.84808, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 169.03397, 321.84808, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 162.71254, 317.2553, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 162.71254, 317.2553, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 157.48415, 311.44858, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 157.48415, 311.44858, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 153.5773, 304.6817, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 153.5773, 304.6817, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 151.16272, 297.25043, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 151.16272, 297.25043, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 150.34598, 289.47952, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 150.34598, 289.47952, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 151.16272, 281.70862, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 151.16272, 281.70862, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 153.5773, 274.27734, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 153.5773, 274.27734, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 157.48415, 267.51047, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 157.48415, 267.51047, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 162.71254, 261.70374, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 162.71254, 261.70374, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 169.03397, 257.11096, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 169.03397, 257.11096, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 176.17215, 253.93283, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 176.17215, 253.93283, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 183.81511, 252.30827, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 183.81511, 252.30827, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 191.62883, 252.30827, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 191.62883, 252.30827, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 199.27179, 253.93283, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 199.27179, 253.93283, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 206.40997, 257.11096, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 206.40997, 257.11096, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 212.7314, 261.70374, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 212.7314, 261.70374, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 217.9598, 267.51047, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 217.9598, 267.51047, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 221.86665, 274.27734, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 221.86665, 274.27734, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 224.28122, 281.70862, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 224.28122, 281.70862, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 225.09798, 289.47952, 1.0, 187.72197, 289.47952, 0.0, 0.0, 0.0, 187.72197, 289.47952, 0.0, 187.72197, 289.47952, 0.0, 1.0, 0.0, 223.13339, 289.85422, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 222.31664, 297.62515, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 222.31664, 297.62515, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 219.90207, 305.05643, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 219.90207, 305.05643, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 215.99521, 311.8233, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 215.99521, 311.8233, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 210.76682, 317.63, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 210.76682, 317.63, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 204.44539, 322.2228, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 204.44539, 322.2228, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 197.3072, 325.4009, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 197.3072, 325.4009, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 189.66425, 327.02548, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 189.66425, 327.02548, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 181.85052, 327.02548, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 181.85052, 327.02548, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 174.20757, 325.4009, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 174.20757, 325.4009, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 167.06938, 322.2228, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 167.06938, 322.2228, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 160.74796, 317.63, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 160.74796, 317.63, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 155.51956, 311.8233, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 155.51956, 311.8233, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 151.61272, 305.05643, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 151.61272, 305.05643, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 149.19815, 297.62515, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 149.19815, 297.62515, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 148.3814, 289.85422, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 148.3814, 289.85422, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 149.19815, 282.0833, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 149.19815, 282.0833, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 151.61272, 274.65204, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 151.61272, 274.65204, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 155.51956, 267.88516, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 155.51956, 267.88516, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 160.74796, 262.07846, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 160.74796, 262.07846, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 167.06938, 257.48566, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 167.06938, 257.48566, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 174.20757, 254.30754, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 174.20757, 254.30754, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 181.85052, 252.68298, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 181.85052, 252.68298, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 189.66425, 252.68298, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 189.66425, 252.68298, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 197.3072, 254.30754, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 197.3072, 254.30754, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 204.44539, 257.48566, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 204.44539, 257.48566, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 210.76682, 262.07846, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 210.76682, 262.07846, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 215.99521, 267.88516, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 215.99521, 267.88516, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 219.90207, 274.65204, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 219.90207, 274.65204, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 222.31664, 282.0833, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 222.31664, 282.0833, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 223.13339, 289.85422, 1.0, 185.75739, 289.85422, 0.0, 0.0, 0.0, 185.75739, 289.85422, 0.0, 185.75739, 289.85422, 0.0, 1.0, 0.0, 221.16971, 290.23367, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 220.35295, 298.00458, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 220.35295, 298.00458, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 217.93839, 305.43585, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 217.93839, 305.43585, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 214.03152, 312.20273, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 214.03152, 312.20273, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 208.80313, 318.00946, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 208.80313, 318.00946, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 202.4817, 322.60223, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 202.4817, 322.60223, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 195.34354, 325.78036, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 195.34354, 325.78036, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 187.70056, 327.40494, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 187.70056, 327.40494, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 179.88686, 327.40494, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 179.88686, 327.40494, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 172.2439, 325.78036, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 172.2439, 325.78036, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 165.10571, 322.60223, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 165.10571, 322.60223, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 158.78429, 318.00946, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 158.78429, 318.00946, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 153.5559, 312.20273, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 153.5559, 312.20273, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 149.64903, 305.43585, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 149.64903, 305.43585, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 147.23447, 298.00458, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 147.23447, 298.00458, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 146.41771, 290.23367, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 146.41771, 290.23367, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 147.23447, 282.46277, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 147.23447, 282.46277, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 149.64903, 275.0315, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 149.64903, 275.0315, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 153.5559, 268.26462, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 153.5559, 268.26462, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 158.78429, 262.4579, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 158.78429, 262.4579, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 165.10571, 257.8651, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 165.10571, 257.8651, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 172.2439, 254.68698, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 172.2439, 254.68698, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 179.88686, 253.06242, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 179.88686, 253.06242, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 187.70056, 253.06242, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 187.70056, 253.06242, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 195.34354, 254.68698, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 195.34354, 254.68698, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 202.4817, 257.8651, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 202.4817, 257.8651, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 208.80313, 262.4579, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 208.80313, 262.4579, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 214.03152, 268.26462, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 214.03152, 268.26462, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 217.93839, 275.0315, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 217.93839, 275.0315, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 220.35295, 282.46277, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 220.35295, 282.46277, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 221.16971, 290.23367, 1.0, 183.79372, 290.23367, 0.0, 0.0, 0.0, 183.79372, 290.23367, 0.0, 183.79372, 290.23367, 0.0, 1.0, 0.0, 219.20695, 290.61786, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 218.3902, 298.38876, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 218.3902, 298.38876, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 215.97563, 305.82004, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 215.97563, 305.82004, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 212.06877, 312.5869, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 212.06877, 312.5869, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 206.84038, 318.39362, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 206.84038, 318.39362, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 200.51895, 322.98642, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 200.51895, 322.98642, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 193.38078, 326.16455, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 193.38078, 326.16455, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 185.73781, 327.7891, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 185.73781, 327.7891, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 177.9241, 327.7891, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 177.9241, 327.7891, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 170.28114, 326.16455, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 170.28114, 326.16455, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 163.14296, 322.98642, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 163.14296, 322.98642, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 156.82153, 318.39362, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 156.82153, 318.39362, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 151.59314, 312.5869, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 151.59314, 312.5869, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 147.68628, 305.82004, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 147.68628, 305.82004, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 145.27171, 298.38876, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 145.27171, 298.38876, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 144.45496, 290.61786, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 144.45496, 290.61786, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 145.27171, 282.84695, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 145.27171, 282.84695, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 147.68628, 275.41565, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 147.68628, 275.41565, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 151.59314, 268.64877, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 151.59314, 268.64877, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 156.82153, 262.84207, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 156.82153, 262.84207, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 163.14296, 258.24927, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 163.14296, 258.24927, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 170.28114, 255.07115, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 170.28114, 255.07115, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 177.9241, 253.4466, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 177.9241, 253.4466, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 185.73781, 253.4466, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 185.73781, 253.4466, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 193.38078, 255.07115, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 193.38078, 255.07115, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 200.51895, 258.24927, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 200.51895, 258.24927, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 206.84038, 262.84207, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 206.84038, 262.84207, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 212.06877, 268.64877, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 212.06877, 268.64877, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 215.97563, 275.41565, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 215.97563, 275.41565, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 218.3902, 282.84695, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 218.3902, 282.84695, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 219.20695, 290.61786, 1.0, 181.83096, 290.61786, 0.0, 0.0, 0.0, 181.83096, 290.61786, 0.0, 181.83096, 290.61786, 0.0, 1.0, 0.0, 217.24513, 291.00674, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 216.42838, 298.77765, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 216.42838, 298.77765, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 214.01381, 306.20895, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 214.01381, 306.20895, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 210.10695, 312.9758, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 210.10695, 312.9758, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 204.87856, 318.78253, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 204.87856, 318.78253, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 198.55713, 323.3753, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 198.55713, 323.3753, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 191.41895, 326.55344, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 191.41895, 326.55344, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 183.77599, 328.178, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 183.77599, 328.178, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 175.96228, 328.178, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 175.96228, 328.178, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 168.31932, 326.55344, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 168.31932, 326.55344, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 161.18114, 323.3753, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 161.18114, 323.3753, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 154.85971, 318.78253, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 154.85971, 318.78253, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 149.63132, 312.9758, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 149.63132, 312.9758, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 145.72446, 306.20895, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 145.72446, 306.20895, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 143.30989, 298.77765, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 143.30989, 298.77765, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 142.49313, 291.00674, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 142.49313, 291.00674, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 143.30989, 283.23584, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 143.30989, 283.23584, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 145.72446, 275.80457, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 145.72446, 275.80457, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 149.63132, 269.0377, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 149.63132, 269.0377, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 154.85971, 263.23096, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 154.85971, 263.23096, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 161.18114, 258.63818, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 161.18114, 258.63818, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 168.31932, 255.46007, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 168.31932, 255.46007, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 175.96228, 253.8355, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 175.96228, 253.8355, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 183.77599, 253.8355, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 183.77599, 253.8355, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 191.41895, 255.46007, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 191.41895, 255.46007, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 198.55713, 258.63818, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 198.55713, 258.63818, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 204.87856, 263.23096, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 204.87856, 263.23096, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 210.10695, 269.0377, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 210.10695, 269.0377, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 214.01381, 275.80457, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 214.01381, 275.80457, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 216.42838, 283.23584, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 216.42838, 283.23584, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 217.24513, 291.00674, 1.0, 179.86914, 291.00674, 0.0, 0.0, 0.0, 179.86914, 291.00674, 0.0, 179.86914, 291.00674, 0.0, 1.0, 0.0, 215.28426, 291.4004, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 214.4675, 299.1713, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 214.4675, 299.1713, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 212.05293, 306.60257, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 212.05293, 306.60257, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 208.14607, 313.36945, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 208.14607, 313.36945, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 202.91768, 319.17615, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 202.91768, 319.17615, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 196.59625, 323.76895, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 196.59625, 323.76895, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 189.45807, 326.94708, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 189.45807, 326.94708, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 181.81511, 328.57162, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 181.81511, 328.57162, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 174.0014, 328.57162, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 174.0014, 328.57162, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 166.35843, 326.94708, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 166.35843, 326.94708, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 159.22025, 323.76895, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 159.22025, 323.76895, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 152.89883, 319.17615, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 152.89883, 319.17615, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 147.67044, 313.36945, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 147.67044, 313.36945, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 143.76358, 306.60257, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 143.76358, 306.60257, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 141.34901, 299.1713, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 141.34901, 299.1713, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 140.53226, 291.4004, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 140.53226, 291.4004, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 141.34901, 283.6295, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 141.34901, 283.6295, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 143.76358, 276.19818, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 143.76358, 276.19818, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 147.67044, 269.4313, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 147.67044, 269.4313, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 152.89883, 263.6246, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 152.89883, 263.6246, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 159.22025, 259.03183, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 159.22025, 259.03183, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 166.35843, 255.8537, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 166.35843, 255.8537, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 174.0014, 254.22913, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 174.0014, 254.22913, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 181.81511, 254.22913, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 181.81511, 254.22913, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 189.45807, 255.8537, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 189.45807, 255.8537, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 196.59625, 259.03183, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 196.59625, 259.03183, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 202.91768, 263.6246, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 202.91768, 263.6246, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 208.14607, 269.4313, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 208.14607, 269.4313, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 212.05293, 276.19818, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 212.05293, 276.19818, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 214.4675, 283.6295, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 214.4675, 283.6295, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 215.28426, 291.4004, 1.0, 177.90825, 291.4004, 0.0, 0.0, 0.0, 177.90825, 291.4004, 0.0, 177.90825, 291.4004, 0.0, 1.0, 0.0, 213.32433, 291.79874, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 212.50757, 299.56964, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 212.50757, 299.56964, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 210.093, 307.00092, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 210.093, 307.00092, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 206.18614, 313.7678, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 206.18614, 313.7678, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 200.95775, 319.57452, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 200.95775, 319.57452, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 194.63632, 324.1673, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 194.63632, 324.1673, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 187.49814, 327.34543, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 187.49814, 327.34543, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 179.85518, 328.97, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 179.85518, 328.97, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 172.04147, 328.97, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 172.04147, 328.97, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 164.39851, 327.34543, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 164.39851, 327.34543, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 157.26033, 324.1673, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 157.26033, 324.1673, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 150.9389, 319.57452, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 150.9389, 319.57452, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 145.71051, 313.7678, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 145.71051, 313.7678, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 141.80365, 307.00092, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 141.80365, 307.00092, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 139.38908, 299.56964, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 139.38908, 299.56964, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 138.57233, 291.79874, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 138.57233, 291.79874, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 139.38908, 284.02783, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 139.38908, 284.02783, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 141.80365, 276.59656, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 141.80365, 276.59656, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 145.71051, 269.82968, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 145.71051, 269.82968, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 150.9389, 264.02295, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 150.9389, 264.02295, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 157.26033, 259.43018, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 157.26033, 259.43018, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 164.39851, 256.25204, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 164.39851, 256.25204, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 172.04147, 254.62749, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 172.04147, 254.62749, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 179.85518, 254.62749, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 179.85518, 254.62749, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 187.49814, 256.25204, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 187.49814, 256.25204, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 194.63632, 259.43018, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 194.63632, 259.43018, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 200.95775, 264.02295, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 200.95775, 264.02295, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 206.18614, 269.82968, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 206.18614, 269.82968, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 210.093, 276.59656, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 210.093, 276.59656, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 212.50757, 284.02783, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 212.50757, 284.02783, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 213.32433, 291.79874, 1.0, 175.94833, 291.79874, 0.0, 0.0, 0.0, 175.94833, 291.79874, 0.0, 175.94833, 291.79874, 0.0, 1.0, 0.0, 211.36537, 292.2018, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 210.54861, 299.97272, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 210.54861, 299.97272, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 208.13403, 307.404, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 208.13403, 307.404, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 204.22719, 314.17087, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 204.22719, 314.17087, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 198.9988, 319.9776, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 198.9988, 319.9776, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 192.67737, 324.57037, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 192.67737, 324.57037, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 185.53918, 327.7485, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 185.53918, 327.7485, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 177.89622, 329.37308, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 177.89622, 329.37308, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 170.0825, 329.37308, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 170.0825, 329.37308, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 162.43954, 327.7485, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 162.43954, 327.7485, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 155.30136, 324.57037, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 155.30136, 324.57037, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 148.97993, 319.9776, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 148.97993, 319.9776, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 143.75154, 314.17087, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 143.75154, 314.17087, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 139.8447, 307.404, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 139.8447, 307.404, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 137.43011, 299.97272, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 137.43011, 299.97272, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 136.61337, 292.2018, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 136.61337, 292.2018, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 137.43011, 284.4309, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 137.43011, 284.4309, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 139.8447, 276.99963, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 139.8447, 276.99963, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 143.75154, 270.23276, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 143.75154, 270.23276, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 148.97993, 264.42603, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 148.97993, 264.42603, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 155.30136, 259.83325, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 155.30136, 259.83325, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 162.43954, 256.65512, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 162.43954, 256.65512, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 170.0825, 255.03056, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 170.0825, 255.03056, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 177.89622, 255.03056, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 177.89622, 255.03056, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 185.53918, 256.65512, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 185.53918, 256.65512, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 192.67737, 259.83325, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 192.67737, 259.83325, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 198.9988, 264.42603, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 198.9988, 264.42603, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 204.22719, 270.23276, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 204.22719, 270.23276, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 208.13403, 276.99963, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 208.13403, 276.99963, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 210.54861, 284.4309, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 210.54861, 284.4309, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 211.36537, 292.2018, 1.0, 173.98936, 292.2018, 0.0, 0.0, 0.0, 173.98936, 292.2018, 0.0, 173.98936, 292.2018, 0.0, 1.0, 0.0, 209.40738, 292.60962, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 208.59062, 300.38052, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 208.59062, 300.38052, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 206.17606, 307.8118, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 206.17606, 307.8118, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 202.2692, 314.57867, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 202.2692, 314.57867, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 197.0408, 320.3854, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 197.0408, 320.3854, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 190.71938, 324.97818, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 190.71938, 324.97818, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 183.5812, 328.1563, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 183.5812, 328.1563, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 175.93823, 329.78085, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 175.93823, 329.78085, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 168.12453, 329.78085, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 168.12453, 329.78085, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 160.48157, 328.1563, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 160.48157, 328.1563, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 153.34338, 324.97818, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 153.34338, 324.97818, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 147.02196, 320.3854, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 147.02196, 320.3854, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 141.79356, 314.57867, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 141.79356, 314.57867, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 137.8867, 307.8118, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 137.8867, 307.8118, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 135.47214, 300.38052, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 135.47214, 300.38052, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 134.65538, 292.60962, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 134.65538, 292.60962, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 135.47214, 284.8387, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 135.47214, 284.8387, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 137.8867, 277.4074, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 137.8867, 277.4074, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 141.79356, 270.64056, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 141.79356, 270.64056, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 147.02196, 264.83383, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 147.02196, 264.83383, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 153.34338, 260.24106, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 153.34338, 260.24106, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 160.48157, 257.06293, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 160.48157, 257.06293, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 168.12453, 255.43835, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 168.12453, 255.43835, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 175.93823, 255.43835, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 175.93823, 255.43835, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 183.5812, 257.06293, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 183.5812, 257.06293, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 190.71938, 260.24106, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 190.71938, 260.24106, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 197.0408, 264.83383, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 197.0408, 264.83383, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 202.2692, 270.64056, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 202.2692, 270.64056, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 206.17606, 277.4074, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 206.17606, 277.4074, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 208.59062, 284.8387, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 208.59062, 284.8387, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 209.40738, 292.60962, 1.0, 172.03139, 292.60962, 0.0, 0.0, 0.0, 172.03139, 292.60962, 0.0, 172.03139, 292.60962, 0.0, 1.0, 0.0, 207.4504, 293.02213, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 206.63364, 300.79303, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 206.63364, 300.79303, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 204.21906, 308.2243, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 204.21906, 308.2243, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 200.31221, 314.99118, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 200.31221, 314.99118, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 195.08382, 320.7979, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 195.08382, 320.7979, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 188.76239, 325.3907, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 188.76239, 325.3907, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 181.6242, 328.56882, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 181.6242, 328.56882, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 173.98125, 330.1934, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 173.98125, 330.1934, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 166.16753, 330.1934, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 166.16753, 330.1934, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 158.52457, 328.56882, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 158.52457, 328.56882, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 151.38638, 325.3907, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 151.38638, 325.3907, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 145.06496, 320.7979, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 145.06496, 320.7979, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 139.83656, 314.99118, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 139.83656, 314.99118, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 135.92972, 308.2243, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 135.92972, 308.2243, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 133.51514, 300.79303, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 133.51514, 300.79303, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 132.6984, 293.02213, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 132.6984, 293.02213, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 133.51514, 285.25122, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 133.51514, 285.25122, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 135.92972, 277.81995, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 135.92972, 277.81995, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 139.83656, 271.05307, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 139.83656, 271.05307, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 145.06496, 265.24634, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 145.06496, 265.24634, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 151.38638, 260.65356, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 151.38638, 260.65356, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 158.52457, 257.47543, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 158.52457, 257.47543, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 166.16753, 255.85088, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 166.16753, 255.85088, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 173.98125, 255.85088, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 173.98125, 255.85088, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 181.6242, 257.47543, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 181.6242, 257.47543, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 188.76239, 260.65356, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 188.76239, 260.65356, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 195.08382, 265.24634, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 195.08382, 265.24634, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 200.31221, 271.05307, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 200.31221, 271.05307, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 204.21906, 277.81995, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 204.21906, 277.81995, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 206.63364, 285.25122, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 206.63364, 285.25122, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 207.4504, 293.02213, 1.0, 170.07439, 293.02213, 0.0, 0.0, 0.0, 170.07439, 293.02213, 0.0, 170.07439, 293.02213, 0.0, 1.0, 0.0, 205.4944, 293.43936, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 204.67764, 301.21027, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 204.67764, 301.21027, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 202.26306, 308.64154, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 202.26306, 308.64154, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 198.35622, 315.40842, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 198.35622, 315.40842, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 193.12782, 321.21515, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 193.12782, 321.21515, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 186.8064, 325.80792, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 186.8064, 325.80792, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 179.66821, 328.98605, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 179.66821, 328.98605, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 172.02525, 330.6106, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 172.02525, 330.6106, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 164.21153, 330.6106, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 164.21153, 330.6106, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 156.56857, 328.98605, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 156.56857, 328.98605, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 149.43039, 325.80792, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 149.43039, 325.80792, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 143.10896, 321.21515, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 143.10896, 321.21515, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 137.88057, 315.40842, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 137.88057, 315.40842, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 133.97372, 308.64154, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 133.97372, 308.64154, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 131.55914, 301.21027, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 131.55914, 301.21027, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 130.74239, 293.43936, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 130.74239, 293.43936, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 131.55914, 285.66846, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 131.55914, 285.66846, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 133.97372, 278.23718, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 133.97372, 278.23718, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 137.88057, 271.4703, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 137.88057, 271.4703, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 143.10896, 265.66357, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 143.10896, 265.66357, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 149.43039, 261.0708, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 149.43039, 261.0708, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 156.56857, 257.89267, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 156.56857, 257.89267, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 164.21153, 256.2681, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 164.21153, 256.2681, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 172.02525, 256.2681, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 172.02525, 256.2681, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 179.66821, 257.89267, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 179.66821, 257.89267, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 186.8064, 261.0708, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 186.8064, 261.0708, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 193.12782, 265.66357, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 193.12782, 265.66357, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 198.35622, 271.4703, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 198.35622, 271.4703, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 202.26306, 278.23718, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 202.26306, 278.23718, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 204.67764, 285.66846, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 204.67764, 285.66846, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 205.4944, 293.43936, 1.0, 168.1184, 293.43936, 0.0, 0.0, 0.0, 168.1184, 293.43936, 0.0, 168.1184, 293.43936, 0.0, 1.0, 0.0, 203.53941, 293.8613, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 202.72266, 301.6322, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 202.72266, 301.6322, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 200.30809, 309.06348, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 200.30809, 309.06348, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 196.40123, 315.83035, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 196.40123, 315.83035, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 191.17284, 321.6371, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 191.17284, 321.6371, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 184.85141, 326.22986, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 184.85141, 326.22986, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 177.71323, 329.408, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 177.71323, 329.408, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 170.07027, 331.03256, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 170.07027, 331.03256, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 162.25655, 331.03256, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 162.25655, 331.03256, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 154.61359, 329.408, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 154.61359, 329.408, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 147.4754, 326.22986, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 147.4754, 326.22986, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 141.15398, 321.6371, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 141.15398, 321.6371, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 135.92558, 315.83035, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 135.92558, 315.83035, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 132.01874, 309.06348, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 132.01874, 309.06348, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 129.60416, 301.6322, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 129.60416, 301.6322, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 128.78741, 293.8613, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 128.78741, 293.8613, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 129.60416, 286.0904, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 129.60416, 286.0904, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 132.01874, 278.65912, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 132.01874, 278.65912, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 135.92558, 271.89224, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 135.92558, 271.89224, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 141.15398, 266.0855, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 141.15398, 266.0855, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 147.4754, 261.49274, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 147.4754, 261.49274, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 154.61359, 258.3146, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 154.61359, 258.3146, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 162.25655, 256.69006, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 162.25655, 256.69006, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 170.07027, 256.69006, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 170.07027, 256.69006, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 177.71323, 258.3146, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 177.71323, 258.3146, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 184.85141, 261.49274, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 184.85141, 261.49274, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 191.17284, 266.0855, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 191.17284, 266.0855, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 196.40123, 271.89224, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 196.40123, 271.89224, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 200.30809, 278.65912, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 200.30809, 278.65912, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 202.72266, 286.0904, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 202.72266, 286.0904, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 203.53941, 293.8613, 1.0, 166.1634, 293.8613, 0.0, 0.0, 0.0, 166.1634, 293.8613, 0.0, 166.1634, 293.8613, 0.0, 1.0, 0.0, 201.58545, 294.28796, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 200.76869, 302.05887, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 200.76869, 302.05887, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 198.35413, 309.49014, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 198.35413, 309.49014, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 194.44727, 316.25702, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 194.44727, 316.25702, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 189.21887, 322.06375, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 189.21887, 322.06375, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 182.89745, 326.65652, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 182.89745, 326.65652, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 175.75926, 329.83466, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 175.75926, 329.83466, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 168.1163, 331.4592, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 168.1163, 331.4592, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 160.3026, 331.4592, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 160.3026, 331.4592, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 152.65962, 329.83466, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 152.65962, 329.83466, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 145.52145, 326.65652, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 145.52145, 326.65652, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 139.20003, 322.06375, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 139.20003, 322.06375, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 133.97163, 316.25702, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 133.97163, 316.25702, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 130.06477, 309.49014, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 130.06477, 309.49014, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 127.6502, 302.05887, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 127.6502, 302.05887, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 126.83345, 294.28796, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 126.83345, 294.28796, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 127.6502, 286.51706, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 127.6502, 286.51706, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 130.06477, 279.08575, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 130.06477, 279.08575, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 133.97163, 272.3189, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 133.97163, 272.3189, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 139.20003, 266.51218, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 139.20003, 266.51218, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 145.52145, 261.9194, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 145.52145, 261.9194, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 152.65962, 258.74127, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 152.65962, 258.74127, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 160.3026, 257.1167, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 160.3026, 257.1167, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 168.1163, 257.1167, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 168.1163, 257.1167, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 175.75926, 258.74127, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 175.75926, 258.74127, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 182.89745, 261.9194, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 182.89745, 261.9194, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 189.21887, 266.51218, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 189.21887, 266.51218, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 194.44727, 272.3189, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 194.44727, 272.3189, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 198.35413, 279.08575, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 198.35413, 279.08575, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 200.76869, 286.51706, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 200.76869, 286.51706, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 201.58545, 294.28796, 1.0, 164.20944, 294.28796, 0.0, 0.0, 0.0, 164.20944, 294.28796, 0.0, 164.20944, 294.28796, 0.0, 1.0, 0.0, 199.63252, 294.71933, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 198.81577, 302.49023, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 198.81577, 302.49023, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 196.4012, 309.9215, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 196.4012, 309.9215, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 192.49434, 316.6884, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 192.49434, 316.6884, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 187.26595, 322.4951, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 187.26595, 322.4951, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 180.94452, 327.0879, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 180.94452, 327.0879, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 173.80634, 330.26602, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 173.80634, 330.26602, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 166.16338, 331.89056, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 166.16338, 331.89056, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 158.34967, 331.89056, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 158.34967, 331.89056, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 150.7067, 330.26602, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 150.7067, 330.26602, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 143.56853, 327.0879, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 143.56853, 327.0879, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 137.2471, 322.4951, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 137.2471, 322.4951, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 132.0187, 316.6884, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 132.0187, 316.6884, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 128.11185, 309.9215, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 128.11185, 309.9215, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 125.69727, 302.49023, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 125.69727, 302.49023, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 124.88052, 294.71933, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 124.88052, 294.71933, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 125.69727, 286.94843, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 125.69727, 286.94843, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 128.11185, 279.51712, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 128.11185, 279.51712, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 132.0187, 272.75024, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 132.0187, 272.75024, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 137.2471, 266.94354, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 137.2471, 266.94354, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 143.56853, 262.35077, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 143.56853, 262.35077, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 150.7067, 259.17264, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 150.7067, 259.17264, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 158.34967, 257.54807, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 158.34967, 257.54807, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 166.16338, 257.54807, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 166.16338, 257.54807, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 173.80634, 259.17264, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 173.80634, 259.17264, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 180.94452, 262.35077, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 180.94452, 262.35077, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 187.26595, 266.94354, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 187.26595, 266.94354, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 192.49434, 272.75024, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 192.49434, 272.75024, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 196.4012, 279.51712, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 196.4012, 279.51712, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 198.81577, 286.94843, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 198.81577, 286.94843, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 199.63252, 294.71933, 1.0, 162.25652, 294.71933, 0.0, 0.0, 0.0, 162.25652, 294.71933, 0.0, 162.25652, 294.71933, 0.0, 1.0, 0.0, 197.68063, 295.1554, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 196.86388, 302.9263, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 196.86388, 302.9263, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 194.44931, 310.35757, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 194.44931, 310.35757, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 190.54247, 317.12445, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 190.54247, 317.12445, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 185.31407, 322.93118, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 185.31407, 322.93118, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 178.99265, 327.52396, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 178.99265, 327.52396, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 171.85446, 330.7021, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 171.85446, 330.7021, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 164.21149, 332.32663, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 164.21149, 332.32663, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 156.39778, 332.32663, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 156.39778, 332.32663, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 148.75482, 330.7021, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 148.75482, 330.7021, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 141.61664, 327.52396, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 141.61664, 327.52396, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 135.29521, 322.93118, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 135.29521, 322.93118, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 130.06682, 317.12445, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 130.06682, 317.12445, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 126.159966, 310.35757, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 126.159966, 310.35757, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 123.74539, 302.9263, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 123.74539, 302.9263, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 122.92864, 295.1554, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 122.92864, 295.1554, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 123.74539, 287.3845, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 123.74539, 287.3845, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 126.159966, 279.9532, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 126.159966, 279.9532, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 130.06682, 273.18634, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 130.06682, 273.18634, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 135.29521, 267.3796, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 135.29521, 267.3796, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 141.61664, 262.78683, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 141.61664, 262.78683, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 148.75482, 259.6087, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 148.75482, 259.6087, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 156.39778, 257.98413, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 156.39778, 257.98413, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 164.21149, 257.98413, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 164.21149, 257.98413, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 171.85446, 259.6087, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 171.85446, 259.6087, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 178.99265, 262.78683, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 178.99265, 262.78683, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 185.31407, 267.3796, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 185.31407, 267.3796, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 190.54247, 273.18634, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 190.54247, 273.18634, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 194.44931, 279.9532, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 194.44931, 279.9532, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 196.86388, 287.3845, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 196.86388, 287.3845, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 197.68063, 295.1554, 1.0, 160.30464, 295.1554, 0.0, 0.0, 0.0, 160.30464, 295.1554, 0.0, 160.30464, 295.1554, 0.0, 1.0, 0.0, 195.72981, 295.59616, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 194.91306, 303.36707, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 194.91306, 303.36707, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 192.49849, 310.79834, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 192.49849, 310.79834, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 188.59163, 317.56522, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 188.59163, 317.56522, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 183.36324, 323.37195, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 183.36324, 323.37195, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 177.04181, 327.96472, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 177.04181, 327.96472, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 169.90363, 331.14285, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 169.90363, 331.14285, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 162.26067, 332.7674, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 162.26067, 332.7674, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 154.44696, 332.7674, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 154.44696, 332.7674, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 146.804, 331.14285, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 146.804, 331.14285, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 139.66582, 327.96472, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 139.66582, 327.96472, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 133.34439, 323.37195, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 133.34439, 323.37195, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 128.116, 317.56522, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 128.116, 317.56522, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 124.20914, 310.79834, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 124.20914, 310.79834, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 121.79457, 303.36707, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 121.79457, 303.36707, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 120.97781, 295.59616, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 120.97781, 295.59616, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 121.79457, 287.82526, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 121.79457, 287.82526, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 124.20914, 280.39398, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 124.20914, 280.39398, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 128.116, 273.6271, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 128.116, 273.6271, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 133.34439, 267.82037, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 133.34439, 267.82037, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 139.66582, 263.2276, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 139.66582, 263.2276, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 146.804, 260.04947, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 146.804, 260.04947, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 154.44696, 258.4249, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 154.44696, 258.4249, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 162.26067, 258.4249, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 162.26067, 258.4249, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 169.90363, 260.04947, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 169.90363, 260.04947, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 177.04181, 263.2276, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 177.04181, 263.2276, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 183.36324, 267.82037, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 183.36324, 267.82037, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 188.59163, 273.6271, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 188.59163, 273.6271, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 192.49849, 280.39398, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 192.49849, 280.39398, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 194.91306, 287.82526, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 194.91306, 287.82526, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 195.72981, 295.59616, 1.0, 158.35382, 295.59616, 0.0, 0.0, 0.0, 158.35382, 295.59616, 0.0, 158.35382, 295.59616, 0.0, 1.0, 0.0, 193.78006, 296.04163, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 192.9633, 303.81253, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 192.9633, 303.81253, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 190.54874, 311.2438, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 190.54874, 311.2438, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 186.64188, 318.01068, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 186.64188, 318.01068, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 181.41348, 323.8174, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 181.41348, 323.8174, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 175.09206, 328.4102, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 175.09206, 328.4102, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 167.95387, 331.58832, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 167.95387, 331.58832, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 160.31091, 333.2129, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 160.31091, 333.2129, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 152.49721, 333.2129, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 152.49721, 333.2129, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 144.85423, 331.58832, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 144.85423, 331.58832, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 137.71605, 328.4102, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 137.71605, 328.4102, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 131.39462, 323.8174, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 131.39462, 323.8174, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 126.16624, 318.01068, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 126.16624, 318.01068, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 122.259384, 311.2438, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 122.259384, 311.2438, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 119.84481, 303.81253, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 119.84481, 303.81253, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 119.02805, 296.04163, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 119.02805, 296.04163, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 119.84481, 288.27072, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 119.84481, 288.27072, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 122.259384, 280.83945, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 122.259384, 280.83945, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 126.16624, 274.07257, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 126.16624, 274.07257, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 131.39462, 268.26584, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 131.39462, 268.26584, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 137.71605, 263.67307, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 137.71605, 263.67307, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 144.85423, 260.49493, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 144.85423, 260.49493, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 152.49721, 258.8704, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 152.49721, 258.8704, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 160.31091, 258.8704, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 160.31091, 258.8704, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 167.95387, 260.49493, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 167.95387, 260.49493, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 175.09206, 263.67307, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 175.09206, 263.67307, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 181.41348, 268.26584, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 181.41348, 268.26584, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 186.64188, 274.07257, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 186.64188, 274.07257, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 190.54874, 280.83945, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 190.54874, 280.83945, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 192.9633, 288.27072, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 192.9633, 288.27072, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 193.78006, 296.04163, 1.0, 156.40405, 296.04163, 0.0, 0.0, 0.0, 156.40405, 296.04163, 0.0, 156.40405, 296.04163, 0.0, 1.0, 0.0, 191.83138, 296.4918, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 191.01462, 304.2627, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 191.01462, 304.2627, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 188.60005, 311.694, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 188.60005, 311.694, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 184.69319, 318.46085, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 184.69319, 318.46085, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 179.4648, 324.26758, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 179.4648, 324.26758, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 173.14337, 328.86035, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 173.14337, 328.86035, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 166.0052, 332.03848, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 166.0052, 332.03848, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 158.36223, 333.66306, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 158.36223, 333.66306, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 150.54852, 333.66306, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 150.54852, 333.66306, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 142.90556, 332.03848, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 142.90556, 332.03848, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 135.76738, 328.86035, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 135.76738, 328.86035, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 129.44595, 324.26758, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 129.44595, 324.26758, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 124.21756, 318.46085, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 124.21756, 318.46085, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 120.3107, 311.694, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 120.3107, 311.694, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 117.89613, 304.2627, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 117.89613, 304.2627, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 117.07938, 296.4918, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 117.07938, 296.4918, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 117.89613, 288.7209, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 117.89613, 288.7209, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 120.3107, 281.2896, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 120.3107, 281.2896, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 124.21756, 274.52274, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 124.21756, 274.52274, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 129.44595, 268.716, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 129.44595, 268.716, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 135.76738, 264.12323, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 135.76738, 264.12323, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 142.90556, 260.9451, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 142.90556, 260.9451, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 150.54852, 259.32056, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 150.54852, 259.32056, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 158.36223, 259.32056, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 158.36223, 259.32056, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 166.0052, 260.9451, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 166.0052, 260.9451, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 173.14337, 264.12323, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 173.14337, 264.12323, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 179.4648, 268.716, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 179.4648, 268.716, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 184.69319, 274.52274, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 184.69319, 274.52274, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 188.60005, 281.2896, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 188.60005, 281.2896, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 191.01462, 288.7209, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 191.01462, 288.7209, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 191.83138, 296.4918, 1.0, 154.45538, 296.4918, 0.0, 0.0, 0.0, 154.45538, 296.4918, 0.0, 154.45538, 296.4918, 0.0, 1.0, 0.0, 189.88379, 296.94666, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 189.06703, 304.71756, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 189.06703, 304.71756, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 186.65247, 312.14886, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 186.65247, 312.14886, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 182.7456, 318.9157, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 182.7456, 318.9157, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 177.51721, 324.72244, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 177.51721, 324.72244, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 171.19579, 329.31522, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 171.19579, 329.31522, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 164.05762, 332.49335, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 164.05762, 332.49335, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 156.41464, 334.11792, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 156.41464, 334.11792, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 148.60094, 334.11792, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 148.60094, 334.11792, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 140.95798, 332.49335, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 140.95798, 332.49335, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 133.8198, 329.31522, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 133.8198, 329.31522, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 127.49837, 324.72244, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 127.49837, 324.72244, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 122.26997, 318.9157, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 122.26997, 318.9157, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 118.36311, 312.14886, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 118.36311, 312.14886, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 115.94855, 304.71756, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 115.94855, 304.71756, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 115.13179, 296.94666, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 115.13179, 296.94666, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 115.94855, 289.17575, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 115.94855, 289.17575, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 118.36311, 281.74448, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 118.36311, 281.74448, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 122.26997, 274.9776, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 122.26997, 274.9776, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 127.49837, 269.17087, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 127.49837, 269.17087, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 133.8198, 264.5781, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 133.8198, 264.5781, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 140.95798, 261.39996, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 140.95798, 261.39996, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 148.60094, 259.77542, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 148.60094, 259.77542, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 156.41464, 259.77542, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 156.41464, 259.77542, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 164.05762, 261.39996, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 164.05762, 261.39996, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 171.19579, 264.5781, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 171.19579, 264.5781, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 177.51721, 269.17087, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 177.51721, 269.17087, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 182.7456, 274.9776, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 182.7456, 274.9776, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 186.65247, 281.74448, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 186.65247, 281.74448, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 189.06703, 289.17575, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 189.06703, 289.17575, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 189.88379, 296.94666, 1.0, 152.5078, 296.94666, 0.0, 0.0, 0.0, 152.5078, 296.94666, 0.0, 152.5078, 296.94666, 0.0, 1.0, 0.0, 187.9373, 297.40622, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 187.12054, 305.17712, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 187.12054, 305.17712, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 184.70598, 312.6084, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 184.70598, 312.6084, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 180.79912, 319.37527, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 180.79912, 319.37527, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 175.57072, 325.182, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 175.57072, 325.182, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 169.2493, 329.77478, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 169.2493, 329.77478, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 162.11113, 332.9529, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 162.11113, 332.9529, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 154.46815, 334.57748, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 154.46815, 334.57748, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 146.65445, 334.57748, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 146.65445, 334.57748, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 139.01149, 332.9529, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 139.01149, 332.9529, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 131.8733, 329.77478, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 131.8733, 329.77478, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 125.55188, 325.182, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 125.55188, 325.182, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 120.32349, 319.37527, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 120.32349, 319.37527, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 116.41663, 312.6084, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 116.41663, 312.6084, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 114.00206, 305.17712, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 114.00206, 305.17712, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 113.1853, 297.40622, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 113.1853, 297.40622, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 114.00206, 289.6353, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 114.00206, 289.6353, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 116.41663, 282.20404, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 116.41663, 282.20404, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 120.32349, 275.43716, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 120.32349, 275.43716, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 125.55188, 269.63043, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 125.55188, 269.63043, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 131.8733, 265.03766, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 131.8733, 265.03766, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 139.01149, 261.85953, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 139.01149, 261.85953, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 146.65445, 260.23495, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 146.65445, 260.23495, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 154.46815, 260.23495, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 154.46815, 260.23495, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 162.11113, 261.85953, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 162.11113, 261.85953, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 169.2493, 265.03766, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 169.2493, 265.03766, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 175.57072, 269.63043, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 175.57072, 269.63043, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 180.79912, 275.43716, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 180.79912, 275.43716, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 184.70598, 282.20404, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 184.70598, 282.20404, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 187.12054, 289.6353, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 187.12054, 289.6353, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 187.9373, 297.40622, 1.0, 150.56131, 297.40622, 0.0, 0.0, 0.0, 150.56131, 297.40622, 0.0, 150.56131, 297.40622, 0.0, 1.0, 0.0, 185.99193, 297.87045, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 185.17517, 305.64136, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 185.17517, 305.64136, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 182.7606, 313.07266, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 182.7606, 313.07266, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 178.85374, 319.83954, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 178.85374, 319.83954, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 173.62535, 325.64624, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 173.62535, 325.64624, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 167.30394, 330.23904, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 167.30394, 330.23904, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 160.16576, 333.41714, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 160.16576, 333.41714, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 152.52278, 335.04172, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 152.52278, 335.04172, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 144.70908, 335.04172, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 144.70908, 335.04172, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 137.06612, 333.41714, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 137.06612, 333.41714, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 129.92793, 330.23904, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 129.92793, 330.23904, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 123.60651, 325.64624, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 123.60651, 325.64624, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 118.37811, 319.83954, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 118.37811, 319.83954, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 114.47126, 313.07266, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 114.47126, 313.07266, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 112.05669, 305.64136, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 112.05669, 305.64136, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 111.23993, 297.87045, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 111.23993, 297.87045, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 112.05669, 290.09955, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 112.05669, 290.09955, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 114.47126, 282.66827, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 114.47126, 282.66827, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 118.37811, 275.9014, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 118.37811, 275.9014, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 123.60651, 270.0947, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 123.60651, 270.0947, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 129.92793, 265.5019, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 129.92793, 265.5019, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 137.06612, 262.3238, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 137.06612, 262.3238, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 144.70908, 260.69922, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 144.70908, 260.69922, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 152.52278, 260.69922, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 152.52278, 260.69922, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 160.16576, 262.3238, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 160.16576, 262.3238, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 167.30394, 265.5019, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 167.30394, 265.5019, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 173.62535, 270.0947, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 173.62535, 270.0947, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 178.85374, 275.9014, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 178.85374, 275.9014, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 182.7606, 282.66827, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 182.7606, 282.66827, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 185.17517, 290.09955, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 185.17517, 290.09955, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 185.99193, 297.87045, 1.0, 148.61594, 297.87045, 0.0, 0.0, 0.0, 148.61594, 297.87045, 0.0, 148.61594, 297.87045, 0.0, 1.0, 0.0, 184.04768, 298.3394, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 183.23093, 306.11032, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 183.23093, 306.11032, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 180.81636, 313.5416, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 180.81636, 313.5416, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 176.9095, 320.30847, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 176.9095, 320.30847, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 171.6811, 326.11517, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 171.6811, 326.11517, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 165.35968, 330.70798, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 165.35968, 330.70798, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 158.2215, 333.88608, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 158.2215, 333.88608, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 150.57854, 335.51065, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 150.57854, 335.51065, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 142.76483, 335.51065, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 142.76483, 335.51065, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 135.12187, 333.88608, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 135.12187, 333.88608, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 127.98369, 330.70798, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 127.98369, 330.70798, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 121.66226, 326.11517, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 121.66226, 326.11517, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 116.43387, 320.30847, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 116.43387, 320.30847, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 112.52701, 313.5416, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 112.52701, 313.5416, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 110.11244, 306.11032, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 110.11244, 306.11032, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 109.295685, 298.3394, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 109.295685, 298.3394, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 110.11244, 290.56848, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 110.11244, 290.56848, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 112.52701, 283.1372, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 112.52701, 283.1372, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 116.43387, 276.37033, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 116.43387, 276.37033, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 121.66226, 270.56363, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 121.66226, 270.56363, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 127.98369, 265.97083, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 127.98369, 265.97083, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 135.12187, 262.79272, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 135.12187, 262.79272, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 142.76483, 261.16815, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 142.76483, 261.16815, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 150.57854, 261.16815, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 150.57854, 261.16815, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 158.2215, 262.79272, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 158.2215, 262.79272, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 165.35968, 265.97083, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 165.35968, 265.97083, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 171.6811, 270.56363, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 171.6811, 270.56363, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 176.9095, 276.37033, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 176.9095, 276.37033, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 180.81636, 283.1372, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 180.81636, 283.1372, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 183.23093, 290.56848, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 183.23093, 290.56848, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 184.04768, 298.3394, 1.0, 146.67169, 298.3394, 0.0, 0.0, 0.0, 146.67169, 298.3394, 0.0, 146.67169, 298.3394, 0.0, 1.0, 0.0, 182.10457, 298.81302, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 181.28781, 306.58392, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 181.28781, 306.58392, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 178.87325, 314.0152, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 178.87325, 314.0152, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 174.96638, 320.78207, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 174.96638, 320.78207, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 169.73799, 326.5888, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 169.73799, 326.5888, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 163.41658, 331.18158, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 163.41658, 331.18158, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 156.2784, 334.3597, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 156.2784, 334.3597, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 148.63542, 335.98425, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 148.63542, 335.98425, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 140.82172, 335.98425, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 140.82172, 335.98425, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 133.17876, 334.3597, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 133.17876, 334.3597, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 126.04057, 331.18158, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 126.04057, 331.18158, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 119.71915, 326.5888, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 119.71915, 326.5888, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 114.49075, 320.78207, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 114.49075, 320.78207, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 110.5839, 314.0152, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 110.5839, 314.0152, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 108.16933, 306.58392, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 108.16933, 306.58392, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 107.35257, 298.81302, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 107.35257, 298.81302, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 108.16933, 291.0421, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 108.16933, 291.0421, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 110.5839, 283.61084, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 110.5839, 283.61084, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 114.49075, 276.84396, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 114.49075, 276.84396, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 119.71915, 271.03723, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 119.71915, 271.03723, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 126.04057, 266.44446, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 126.04057, 266.44446, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 133.17876, 263.26633, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 133.17876, 263.26633, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 140.82172, 261.64175, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 140.82172, 261.64175, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 148.63542, 261.64175, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 148.63542, 261.64175, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 156.2784, 263.26633, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 156.2784, 263.26633, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 163.41658, 266.44446, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 163.41658, 266.44446, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 169.73799, 271.03723, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 169.73799, 271.03723, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 174.96638, 276.84396, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 174.96638, 276.84396, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 178.87325, 283.61084, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 178.87325, 283.61084, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 181.28781, 291.0421, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 181.28781, 291.0421, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 182.10457, 298.81302, 1.0, 144.72858, 298.81302, 0.0, 0.0, 0.0, 144.72858, 298.81302, 0.0, 144.72858, 298.81302, 0.0, 1.0, 0.0, 180.16261, 299.29132, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 179.34586, 307.06223, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 179.34586, 307.06223, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 176.93129, 314.4935, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 176.93129, 314.4935, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 173.02443, 321.26038, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 173.02443, 321.26038, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 167.79604, 327.0671, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 167.79604, 327.0671, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 161.47461, 331.65988, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 161.47461, 331.65988, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 154.33643, 334.838, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 154.33643, 334.838, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 146.69347, 336.46255, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 146.69347, 336.46255, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 138.87975, 336.46255, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 138.87975, 336.46255, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 131.23679, 334.838, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 131.23679, 334.838, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 124.09861, 331.65988, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 124.09861, 331.65988, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 117.77718, 327.0671, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 117.77718, 327.0671, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 112.54879, 321.26038, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 112.54879, 321.26038, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 108.64193, 314.4935, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 108.64193, 314.4935, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 106.22736, 307.06223, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 106.22736, 307.06223, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 105.41061, 299.29132, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 105.41061, 299.29132, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 106.22736, 291.52042, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 106.22736, 291.52042, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 108.64193, 284.08914, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 108.64193, 284.08914, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 112.54879, 277.32227, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 112.54879, 277.32227, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 117.77718, 271.51553, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 117.77718, 271.51553, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 124.09861, 266.92276, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 124.09861, 266.92276, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 131.23679, 263.74463, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 131.23679, 263.74463, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 138.87975, 262.12006, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 138.87975, 262.12006, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 146.69347, 262.12006, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 146.69347, 262.12006, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 154.33643, 263.74463, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 154.33643, 263.74463, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 161.47461, 266.92276, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 161.47461, 266.92276, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 167.79604, 271.51553, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 167.79604, 271.51553, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 173.02443, 277.32227, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 173.02443, 277.32227, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 176.93129, 284.08914, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 176.93129, 284.08914, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 179.34586, 291.52042, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 179.34586, 291.52042, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 180.16261, 299.29132, 1.0, 142.7866, 299.29132, 0.0, 0.0, 0.0, 142.7866, 299.29132, 0.0, 142.7866, 299.29132, 0.0, 1.0, 0.0, 178.2218, 299.7743, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 177.40504, 307.5452, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 177.40504, 307.5452, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 174.99048, 314.97647, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 174.99048, 314.97647, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 171.08362, 321.74335, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 171.08362, 321.74335, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 165.85522, 327.55008, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 165.85522, 327.55008, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 159.5338, 332.14285, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 159.5338, 332.14285, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 152.39561, 335.32098, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 152.39561, 335.32098, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 144.75266, 336.94556, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 144.75266, 336.94556, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 136.93895, 336.94556, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 136.93895, 336.94556, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 129.29599, 335.32098, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 129.29599, 335.32098, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 122.1578, 332.14285, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 122.1578, 332.14285, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 115.83638, 327.55008, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 115.83638, 327.55008, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 110.60799, 321.74335, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 110.60799, 321.74335, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 106.701126, 314.97647, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 106.701126, 314.97647, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 104.28656, 307.5452, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 104.28656, 307.5452, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 103.4698, 299.7743, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 103.4698, 299.7743, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 104.28656, 292.0034, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 104.28656, 292.0034, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 106.701126, 284.5721, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 106.701126, 284.5721, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 110.60799, 277.80524, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 110.60799, 277.80524, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 115.83638, 271.9985, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 115.83638, 271.9985, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 122.1578, 267.40573, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 122.1578, 267.40573, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 129.29599, 264.2276, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 129.29599, 264.2276, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 136.93895, 262.60306, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 136.93895, 262.60306, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 144.75266, 262.60306, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 144.75266, 262.60306, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 152.39561, 264.2276, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 152.39561, 264.2276, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 159.5338, 267.40573, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 159.5338, 267.40573, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 165.85522, 271.9985, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 165.85522, 271.9985, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 171.08362, 277.80524, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 171.08362, 277.80524, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 174.99048, 284.5721, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 174.99048, 284.5721, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 177.40504, 292.0034, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 177.40504, 292.0034, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 178.2218, 299.7743, 1.0, 140.8458, 299.7743, 0.0, 0.0, 0.0, 140.8458, 299.7743, 0.0, 140.8458, 299.7743, 0.0, 1.0, 0.0, 176.28217, 300.26196, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 175.46541, 308.03287, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 175.46541, 308.03287, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 173.05084, 315.46414, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 173.05084, 315.46414, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 169.14398, 322.23102, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 169.14398, 322.23102, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 163.91559, 328.03772, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 163.91559, 328.03772, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 157.59416, 332.63052, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 157.59416, 332.63052, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 150.45598, 335.80862, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 150.45598, 335.80862, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 142.81302, 337.4332, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 142.81302, 337.4332, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 134.99931, 337.4332, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 134.99931, 337.4332, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 127.356346, 335.80862, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 127.356346, 335.80862, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 120.21816, 332.63052, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 120.21816, 332.63052, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 113.896736, 328.03772, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 113.896736, 328.03772, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 108.66834, 322.23102, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 108.66834, 322.23102, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 104.76149, 315.46414, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 104.76149, 315.46414, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 102.346924, 308.03287, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 102.346924, 308.03287, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 101.53017, 300.26196, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 101.53017, 300.26196, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 102.346924, 292.49106, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 102.346924, 292.49106, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 104.76149, 285.05975, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 104.76149, 285.05975, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 108.66834, 278.29288, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 108.66834, 278.29288, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 113.896736, 272.48618, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 113.896736, 272.48618, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 120.21816, 267.89337, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 120.21816, 267.89337, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 127.356346, 264.71527, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 127.356346, 264.71527, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 134.99931, 263.0907, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 134.99931, 263.0907, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 142.81302, 263.0907, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 142.81302, 263.0907, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 150.45598, 264.71527, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 150.45598, 264.71527, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 157.59416, 267.89337, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 157.59416, 267.89337, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 163.91559, 272.48618, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 163.91559, 272.48618, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 169.14398, 278.29288, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 169.14398, 278.29288, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 173.05084, 285.05975, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 173.05084, 285.05975, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 175.46541, 292.49106, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 175.46541, 292.49106, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 176.28217, 300.26196, 1.0, 138.90616, 300.26196, 0.0, 0.0, 0.0, 138.90616, 300.26196, 0.0, 138.90616, 300.26196, 0.0, 1.0, 0.0, 174.3437, 300.75427, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 173.52695, 308.52518, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 173.52695, 308.52518, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 171.11238, 315.95648, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 171.11238, 315.95648, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 167.20554, 322.72333, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 167.20554, 322.72333, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 161.97714, 328.53006, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 161.97714, 328.53006, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 155.65572, 333.12283, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 155.65572, 333.12283, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 148.51753, 336.30096, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 148.51753, 336.30096, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 140.87457, 337.92554, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 140.87457, 337.92554, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 133.06085, 337.92554, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 133.06085, 337.92554, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 125.41789, 336.30096, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 125.41789, 336.30096, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 118.27971, 333.12283, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 118.27971, 333.12283, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 111.95828, 328.53006, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 111.95828, 328.53006, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 106.72989, 322.72333, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 106.72989, 322.72333, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 102.82304, 315.95648, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 102.82304, 315.95648, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 100.40846, 308.52518, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 100.40846, 308.52518, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 99.59171, 300.75427, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 99.59171, 300.75427, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 100.40846, 292.98337, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 100.40846, 292.98337, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 102.82304, 285.5521, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 102.82304, 285.5521, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 106.72989, 278.78522, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 106.72989, 278.78522, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 111.95828, 272.9785, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 111.95828, 272.9785, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 118.27971, 268.3857, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 118.27971, 268.3857, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 125.41789, 265.20758, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 125.41789, 265.20758, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 133.06085, 263.58304, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 133.06085, 263.58304, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 140.87457, 263.58304, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 140.87457, 263.58304, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 148.51753, 265.20758, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 148.51753, 265.20758, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 155.65572, 268.3857, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 155.65572, 268.3857, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 161.97714, 272.9785, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 161.97714, 272.9785, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 167.20554, 278.78522, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 167.20554, 278.78522, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 171.11238, 285.5521, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 171.11238, 285.5521, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 173.52695, 292.98337, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 173.52695, 292.98337, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 174.3437, 300.75427, 1.0, 136.96771, 300.75427, 0.0, 0.0, 0.0, 136.96771, 300.75427, 0.0, 136.96771, 300.75427, 0.0, 1.0, 0.0, 172.40645, 301.25128, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 171.58969, 309.0222, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 171.58969, 309.0222, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 169.17513, 316.45346, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 169.17513, 316.45346, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 165.26826, 323.22034, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 165.26826, 323.22034, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 160.03987, 329.02707, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 160.03987, 329.02707, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 153.71844, 333.61984, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 153.71844, 333.61984, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 146.58026, 336.79797, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 146.58026, 336.79797, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 138.9373, 338.42252, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 138.9373, 338.42252, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 131.1236, 338.42252, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 131.1236, 338.42252, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 123.48063, 336.79797, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 123.48063, 336.79797, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 116.342445, 333.61984, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 116.342445, 333.61984, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 110.02102, 329.02707, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 110.02102, 329.02707, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 104.792625, 323.22034, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 104.792625, 323.22034, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 100.88577, 316.45346, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 100.88577, 316.45346, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 98.4712, 309.0222, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 98.4712, 309.0222, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 97.65445, 301.25128, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 97.65445, 301.25128, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 98.4712, 293.48038, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 98.4712, 293.48038, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 100.88577, 286.0491, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 100.88577, 286.0491, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 104.792625, 279.28223, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 104.792625, 279.28223, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 110.02102, 273.4755, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 110.02102, 273.4755, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 116.342445, 268.88272, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 116.342445, 268.88272, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 123.48063, 265.7046, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 123.48063, 265.7046, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 131.1236, 264.08002, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 131.1236, 264.08002, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 138.9373, 264.08002, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 138.9373, 264.08002, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 146.58026, 265.7046, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 146.58026, 265.7046, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 153.71844, 268.88272, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 153.71844, 268.88272, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 160.03987, 273.4755, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 160.03987, 273.4755, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 165.26826, 279.28223, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 165.26826, 279.28223, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 169.17513, 286.0491, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 169.17513, 286.0491, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 171.58969, 293.48038, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 171.58969, 293.48038, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 172.40645, 301.25128, 1.0, 135.03044, 301.25128, 0.0, 0.0, 0.0, 135.03044, 301.25128, 0.0, 135.03044, 301.25128, 0.0, 1.0, 0.0, 170.47038, 301.75293, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 169.65363, 309.52386, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 169.65363, 309.52386, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 167.23906, 316.95514, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 167.23906, 316.95514, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 163.3322, 323.72202, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 163.3322, 323.72202, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 158.1038, 329.52872, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 158.1038, 329.52872, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 151.78238, 334.12152, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 151.78238, 334.12152, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 144.64421, 337.29962, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 144.64421, 337.29962, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 137.00124, 338.9242, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 137.00124, 338.9242, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 129.18753, 338.9242, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 129.18753, 338.9242, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 121.54456, 337.29962, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 121.54456, 337.29962, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 114.40639, 334.12152, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 114.40639, 334.12152, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 108.08496, 329.52872, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 108.08496, 329.52872, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 102.85657, 323.72202, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 102.85657, 323.72202, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 98.94971, 316.95514, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 98.94971, 316.95514, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 96.53514, 309.52386, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 96.53514, 309.52386, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 95.71838, 301.75293, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 95.71838, 301.75293, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 96.53514, 293.98203, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 96.53514, 293.98203, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 98.94971, 286.55075, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 98.94971, 286.55075, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 102.85657, 279.78387, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 102.85657, 279.78387, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 108.08496, 273.97717, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 108.08496, 273.97717, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 114.40639, 269.38437, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 114.40639, 269.38437, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 121.54456, 266.20627, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 121.54456, 266.20627, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 129.18753, 264.5817, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 129.18753, 264.5817, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 137.00124, 264.5817, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 137.00124, 264.5817, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 144.64421, 266.20627, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 144.64421, 266.20627, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 151.78238, 269.38437, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 151.78238, 269.38437, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 158.1038, 273.97717, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 158.1038, 273.97717, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 163.3322, 279.78387, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 163.3322, 279.78387, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 167.23906, 286.55075, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 167.23906, 286.55075, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 169.65363, 293.98203, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 169.65363, 293.98203, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 170.47038, 301.75293, 1.0, 133.09439, 301.75293, 0.0, 0.0, 0.0, 133.09439, 301.75293, 0.0, 133.09439, 301.75293, 0.0, 1.0, 0.0, 168.53554, 302.25928, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 167.71878, 310.03018, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 167.71878, 310.03018, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 165.30421, 317.46146, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 165.30421, 317.46146, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 161.39735, 324.22833, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 161.39735, 324.22833, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 156.16896, 330.03506, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 156.16896, 330.03506, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 149.84753, 334.62784, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 149.84753, 334.62784, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 142.70937, 337.80597, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 142.70937, 337.80597, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 135.06639, 339.4305, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 135.06639, 339.4305, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 127.252686, 339.4305, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 127.252686, 339.4305, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 119.60972, 337.80597, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 119.60972, 337.80597, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 112.47154, 334.62784, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 112.47154, 334.62784, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 106.150116, 330.03506, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 106.150116, 330.03506, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 100.92172, 324.22833, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 100.92172, 324.22833, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 97.01486, 317.46146, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 97.01486, 317.46146, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 94.600296, 310.03018, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 94.600296, 310.03018, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 93.78354, 302.25928, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 93.78354, 302.25928, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 94.600296, 294.48837, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 94.600296, 294.48837, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 97.01486, 287.0571, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 97.01486, 287.0571, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 100.92172, 280.29022, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 100.92172, 280.29022, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 106.150116, 274.4835, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 106.150116, 274.4835, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 112.47154, 269.89072, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 112.47154, 269.89072, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 119.60972, 266.7126, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 119.60972, 266.7126, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 127.252686, 265.088, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 127.252686, 265.088, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 135.06639, 265.088, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 135.06639, 265.088, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 142.70937, 266.7126, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 142.70937, 266.7126, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 149.84753, 269.89072, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 149.84753, 269.89072, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 156.16896, 274.4835, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 156.16896, 274.4835, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 161.39735, 280.29022, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 161.39735, 280.29022, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 165.30421, 287.0571, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 165.30421, 287.0571, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 167.71878, 294.48837, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 167.71878, 294.48837, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 168.53554, 302.25928, 1.0, 131.15955, 302.25928, 0.0, 0.0, 0.0, 131.15955, 302.25928, 0.0, 131.15955, 302.25928, 0.0, 1.0, 0.0, 166.60191, 302.77026, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 165.78517, 310.54117, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 165.78517, 310.54117, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 163.37059, 317.97244, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 163.37059, 317.97244, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 159.46375, 324.73932, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 159.46375, 324.73932, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 154.23535, 330.54605, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 154.23535, 330.54605, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 147.91393, 335.13882, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 147.91393, 335.13882, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 140.77574, 338.31696, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 140.77574, 338.31696, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 133.13278, 339.94153, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 133.13278, 339.94153, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 125.31906, 339.94153, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 125.31906, 339.94153, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 117.6761, 338.31696, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 117.6761, 338.31696, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 110.53792, 335.13882, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 110.53792, 335.13882, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 104.21649, 330.54605, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 104.21649, 330.54605, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 98.9881, 324.73932, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 98.9881, 324.73932, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 95.081245, 317.97244, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 95.081245, 317.97244, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 92.66668, 310.54117, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 92.66668, 310.54117, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 91.84992, 302.77026, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 91.84992, 302.77026, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 92.66668, 294.99936, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 92.66668, 294.99936, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 95.081245, 287.56808, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 95.081245, 287.56808, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 98.9881, 280.8012, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 98.9881, 280.8012, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 104.21649, 274.99448, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 104.21649, 274.99448, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 110.53792, 270.4017, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 110.53792, 270.4017, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 117.6761, 267.22357, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 117.6761, 267.22357, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 125.31906, 265.59903, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 125.31906, 265.59903, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 133.13278, 265.59903, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 133.13278, 265.59903, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 140.77574, 267.22357, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 140.77574, 267.22357, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 147.91393, 270.4017, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 147.91393, 270.4017, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 154.23535, 274.99448, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 154.23535, 274.99448, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 159.46375, 280.8012, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 159.46375, 280.8012, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 163.37059, 287.56808, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 163.37059, 287.56808, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 165.78517, 294.99936, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 165.78517, 294.99936, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 166.60191, 302.77026, 1.0, 129.22592, 302.77026, 0.0, 0.0, 0.0, 129.22592, 302.77026, 0.0, 129.22592, 302.77026, 0.0, 1.0, 0.0, 164.66954, 303.28592, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 163.85278, 311.05682, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 163.85278, 311.05682, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 161.43822, 318.4881, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 161.43822, 318.4881, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 157.53136, 325.25497, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 157.53136, 325.25497, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 152.30296, 331.0617, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 152.30296, 331.0617, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 145.98154, 335.65448, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 145.98154, 335.65448, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 138.84335, 338.8326, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 138.84335, 338.8326, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 131.2004, 340.45715, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 131.2004, 340.45715, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 123.38668, 340.45715, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 123.38668, 340.45715, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 115.74372, 338.8326, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 115.74372, 338.8326, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 108.60554, 335.65448, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 108.60554, 335.65448, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 102.28411, 331.0617, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 102.28411, 331.0617, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 97.05572, 325.25497, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 97.05572, 325.25497, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 93.148865, 318.4881, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 93.148865, 318.4881, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 90.73429, 311.05682, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 90.73429, 311.05682, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 89.91754, 303.28592, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 89.91754, 303.28592, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 90.73429, 295.515, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 90.73429, 295.515, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 93.148865, 288.08374, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 93.148865, 288.08374, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 97.05572, 281.31686, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 97.05572, 281.31686, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 102.28411, 275.51013, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 102.28411, 275.51013, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 108.60554, 270.91736, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 108.60554, 270.91736, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 115.74372, 267.73923, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 115.74372, 267.73923, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 123.38668, 266.11465, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 123.38668, 266.11465, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 131.2004, 266.11465, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 131.2004, 266.11465, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 138.84335, 267.73923, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 138.84335, 267.73923, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 145.98154, 270.91736, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 145.98154, 270.91736, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 152.30296, 275.51013, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 152.30296, 275.51013, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 157.53136, 281.31686, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 157.53136, 281.31686, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 161.43822, 288.08374, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 161.43822, 288.08374, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 163.85278, 295.515, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 163.85278, 295.515, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 164.66954, 303.28592, 1.0, 127.29354, 303.28592, 0.0, 0.0, 0.0, 127.29354, 303.28592, 0.0, 127.29354, 303.28592, 0.0, 1.0, 0.0, 162.7384, 303.8062, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 161.92165, 311.57712, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 161.92165, 311.57712, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 159.50708, 319.00842, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 159.50708, 319.00842, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 155.60022, 325.7753, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 155.60022, 325.7753, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 150.37183, 331.582, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 150.37183, 331.582, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 144.0504, 336.1748, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 144.0504, 336.1748, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 136.91222, 339.3529, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 136.91222, 339.3529, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 129.26926, 340.97748, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 129.26926, 340.97748, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 121.45555, 340.97748, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 121.45555, 340.97748, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 113.812584, 339.3529, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 113.812584, 339.3529, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 106.6744, 336.1748, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 106.6744, 336.1748, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 100.35298, 331.582, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 100.35298, 331.582, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 95.12459, 325.7753, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 95.12459, 325.7753, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 91.21773, 319.00842, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 91.21773, 319.00842, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 88.80316, 311.57712, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 88.80316, 311.57712, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 87.986404, 303.8062, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 87.986404, 303.8062, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 88.80316, 296.0353, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 88.80316, 296.0353, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 91.21773, 288.60403, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 91.21773, 288.60403, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 95.12459, 281.83716, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 95.12459, 281.83716, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 100.35298, 276.03046, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 100.35298, 276.03046, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 106.6744, 271.43765, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 106.6744, 271.43765, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 113.812584, 268.25955, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 113.812584, 268.25955, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 121.45555, 266.63498, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 121.45555, 266.63498, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 129.26926, 266.63498, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 129.26926, 266.63498, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 136.91222, 268.25955, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 136.91222, 268.25955, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 144.0504, 271.43765, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 144.0504, 271.43765, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 150.37183, 276.03046, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 150.37183, 276.03046, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 155.60022, 281.83716, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 155.60022, 281.83716, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 159.50708, 288.60403, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 159.50708, 288.60403, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 161.92165, 296.0353, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0, 161.92165, 296.0353, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 162.7384, 303.8062, 1.0, 125.362404, 303.8062, 0.0, 0.0, 0.0, 125.362404, 303.8062, 0.0, 125.362404, 303.8062, 0.0, 1.0, 0.0
	]

)
