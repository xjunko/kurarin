module tinyfiledialogs

// Public
pub fn open_file_picker(title string, starting_path string, filters []string, filters_name string, multiple bool) string {
	return ''
}
